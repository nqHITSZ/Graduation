`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/10/11 13:25:03
// Design Name: 
// Module Name: buffer52
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//NOTE: The filter center is reg_26_26; reg_26_26 represent (27,27) (start at 1 not 0)
module  window52 
#(
    parameter DATA_WIDTH = 28,
    parameter IMAGE_WIDTH = 640,
    parameter REGSNUM = 52
)
(
    input wire [DATA_WIDTH - 1:0]  din,
    input wire din_valid,
    input wire clk,
    input wire rst,
    
//    input [9:0] i_row_cnt, i_col_cnt,
//    output [9:0] o_row_cnt, o_col_cnt,
    
    output wire  dout_valid,
    //output format:reg_x_y
    output wire [DATA_WIDTH - 1:0] reg_10_01,
    output wire [DATA_WIDTH - 1:0] reg_43_01,
    output wire [DATA_WIDTH - 1:0] reg_12_04,
    output wire [DATA_WIDTH - 1:0] reg_41_04,
    output wire [DATA_WIDTH - 1:0] reg_14_07,
    output wire [DATA_WIDTH - 1:0] reg_39_07,
    output wire [DATA_WIDTH - 1:0] reg_09_09,
    output wire [DATA_WIDTH - 1:0] reg_26_09,
    output wire [DATA_WIDTH - 1:0] reg_27_09,
    output wire [DATA_WIDTH - 1:0] reg_44_09,
    output wire [DATA_WIDTH - 1:0] reg_01_10,
    output wire [DATA_WIDTH - 1:0] reg_16_10,
    output wire [DATA_WIDTH - 1:0] reg_18_10,
    output wire [DATA_WIDTH - 1:0] reg_35_10,
    output wire [DATA_WIDTH - 1:0] reg_37_10,
    output wire [DATA_WIDTH - 1:0] reg_52_10,
    output wire [DATA_WIDTH - 1:0] reg_11_11,
    output wire [DATA_WIDTH - 1:0] reg_26_11,
    output wire [DATA_WIDTH - 1:0] reg_27_11,
    output wire [DATA_WIDTH - 1:0] reg_42_11,
    output wire [DATA_WIDTH - 1:0] reg_04_12,
    output wire [DATA_WIDTH - 1:0] reg_19_12,
    output wire [DATA_WIDTH - 1:0] reg_34_12,
    output wire [DATA_WIDTH - 1:0] reg_49_12,
    output wire [DATA_WIDTH - 1:0] reg_13_13,
    output wire [DATA_WIDTH - 1:0] reg_18_13,
    output wire [DATA_WIDTH - 1:0] reg_26_13,
    output wire [DATA_WIDTH - 1:0] reg_27_13,
    output wire [DATA_WIDTH - 1:0] reg_35_13,
    output wire [DATA_WIDTH - 1:0] reg_40_13,
    output wire [DATA_WIDTH - 1:0] reg_07_14,
    output wire [DATA_WIDTH - 1:0] reg_20_14,
    output wire [DATA_WIDTH - 1:0] reg_33_14,
    output wire [DATA_WIDTH - 1:0] reg_46_14,
    output wire [DATA_WIDTH - 1:0] reg_15_15,
    output wire [DATA_WIDTH - 1:0] reg_26_15,
    output wire [DATA_WIDTH - 1:0] reg_27_15,
    output wire [DATA_WIDTH - 1:0] reg_38_15,
    output wire [DATA_WIDTH - 1:0] reg_10_16,
    output wire [DATA_WIDTH - 1:0] reg_20_16,
    output wire [DATA_WIDTH - 1:0] reg_21_16,
    output wire [DATA_WIDTH - 1:0] reg_32_16,
    output wire [DATA_WIDTH - 1:0] reg_33_16,
    output wire [DATA_WIDTH - 1:0] reg_43_16,
    output wire [DATA_WIDTH - 1:0] reg_17_17,
    output wire [DATA_WIDTH - 1:0] reg_26_17,
    output wire [DATA_WIDTH - 1:0] reg_27_17,
    output wire [DATA_WIDTH - 1:0] reg_36_17,
    output wire [DATA_WIDTH - 1:0] reg_10_18,
    output wire [DATA_WIDTH - 1:0] reg_13_18,
    output wire [DATA_WIDTH - 1:0] reg_22_18,
    output wire [DATA_WIDTH - 1:0] reg_31_18,
    output wire [DATA_WIDTH - 1:0] reg_40_18,
    output wire [DATA_WIDTH - 1:0] reg_43_18,
    output wire [DATA_WIDTH - 1:0] reg_12_19,
    output wire [DATA_WIDTH - 1:0] reg_19_19,
    output wire [DATA_WIDTH - 1:0] reg_22_19,
    output wire [DATA_WIDTH - 1:0] reg_26_19,
    output wire [DATA_WIDTH - 1:0] reg_27_19,
    output wire [DATA_WIDTH - 1:0] reg_31_19,
    output wire [DATA_WIDTH - 1:0] reg_34_19,
    output wire [DATA_WIDTH - 1:0] reg_41_19,
    output wire [DATA_WIDTH - 1:0] reg_14_20,
    output wire [DATA_WIDTH - 1:0] reg_16_20,
    output wire [DATA_WIDTH - 1:0] reg_23_20,
    output wire [DATA_WIDTH - 1:0] reg_30_20,
    output wire [DATA_WIDTH - 1:0] reg_37_20,
    output wire [DATA_WIDTH - 1:0] reg_39_20,
    output wire [DATA_WIDTH - 1:0] reg_16_21,
    output wire [DATA_WIDTH - 1:0] reg_21_21,
    output wire [DATA_WIDTH - 1:0] reg_26_21,
    output wire [DATA_WIDTH - 1:0] reg_27_21,
    output wire [DATA_WIDTH - 1:0] reg_32_21,
    output wire [DATA_WIDTH - 1:0] reg_37_21,
    output wire [DATA_WIDTH - 1:0] reg_18_22,
    output wire [DATA_WIDTH - 1:0] reg_19_22,
    output wire [DATA_WIDTH - 1:0] reg_24_22,
    output wire [DATA_WIDTH - 1:0] reg_29_22,
    output wire [DATA_WIDTH - 1:0] reg_34_22,
    output wire [DATA_WIDTH - 1:0] reg_35_22,
    output wire [DATA_WIDTH - 1:0] reg_20_23,
    output wire [DATA_WIDTH - 1:0] reg_23_23,
    output wire [DATA_WIDTH - 1:0] reg_26_23,
    output wire [DATA_WIDTH - 1:0] reg_27_23,
    output wire [DATA_WIDTH - 1:0] reg_30_23,
    output wire [DATA_WIDTH - 1:0] reg_33_23,
    output wire [DATA_WIDTH - 1:0] reg_22_24,
    output wire [DATA_WIDTH - 1:0] reg_25_24,
    output wire [DATA_WIDTH - 1:0] reg_28_24,
    output wire [DATA_WIDTH - 1:0] reg_31_24,
    output wire [DATA_WIDTH - 1:0] reg_24_25,
    output wire [DATA_WIDTH - 1:0] reg_29_25,
    output wire [DATA_WIDTH - 1:0] reg_09_26,
    output wire [DATA_WIDTH - 1:0] reg_11_26,
    output wire [DATA_WIDTH - 1:0] reg_13_26,
    output wire [DATA_WIDTH - 1:0] reg_15_26,
    output wire [DATA_WIDTH - 1:0] reg_17_26,
    output wire [DATA_WIDTH - 1:0] reg_19_26,
    output wire [DATA_WIDTH - 1:0] reg_21_26,
    output wire [DATA_WIDTH - 1:0] reg_23_26,
    output wire [DATA_WIDTH - 1:0] reg_26_26,
    output wire [DATA_WIDTH - 1:0] reg_27_26,
    output wire [DATA_WIDTH - 1:0] reg_30_26,
    output wire [DATA_WIDTH - 1:0] reg_32_26,
    output wire [DATA_WIDTH - 1:0] reg_34_26,
    output wire [DATA_WIDTH - 1:0] reg_36_26,
    output wire [DATA_WIDTH - 1:0] reg_38_26,
    output wire [DATA_WIDTH - 1:0] reg_40_26,
    output wire [DATA_WIDTH - 1:0] reg_42_26,
    output wire [DATA_WIDTH - 1:0] reg_44_26,
    output wire [DATA_WIDTH - 1:0] reg_09_27,
    output wire [DATA_WIDTH - 1:0] reg_11_27,
    output wire [DATA_WIDTH - 1:0] reg_13_27,
    output wire [DATA_WIDTH - 1:0] reg_15_27,
    output wire [DATA_WIDTH - 1:0] reg_17_27,
    output wire [DATA_WIDTH - 1:0] reg_19_27,
    output wire [DATA_WIDTH - 1:0] reg_21_27,
    output wire [DATA_WIDTH - 1:0] reg_23_27,
    output wire [DATA_WIDTH - 1:0] reg_26_27,
    output wire [DATA_WIDTH - 1:0] reg_27_27,
    output wire [DATA_WIDTH - 1:0] reg_30_27,
    output wire [DATA_WIDTH - 1:0] reg_32_27,
    output wire [DATA_WIDTH - 1:0] reg_34_27,
    output wire [DATA_WIDTH - 1:0] reg_36_27,
    output wire [DATA_WIDTH - 1:0] reg_38_27,
    output wire [DATA_WIDTH - 1:0] reg_40_27,
    output wire [DATA_WIDTH - 1:0] reg_42_27,
    output wire [DATA_WIDTH - 1:0] reg_44_27,
    output wire [DATA_WIDTH - 1:0] reg_24_28,
    output wire [DATA_WIDTH - 1:0] reg_29_28,
    output wire [DATA_WIDTH - 1:0] reg_22_29,
    output wire [DATA_WIDTH - 1:0] reg_25_29,
    output wire [DATA_WIDTH - 1:0] reg_28_29,
    output wire [DATA_WIDTH - 1:0] reg_31_29,
    output wire [DATA_WIDTH - 1:0] reg_20_30,
    output wire [DATA_WIDTH - 1:0] reg_23_30,
    output wire [DATA_WIDTH - 1:0] reg_26_30,
    output wire [DATA_WIDTH - 1:0] reg_27_30,
    output wire [DATA_WIDTH - 1:0] reg_30_30,
    output wire [DATA_WIDTH - 1:0] reg_33_30,
    output wire [DATA_WIDTH - 1:0] reg_18_31,
    output wire [DATA_WIDTH - 1:0] reg_19_31,
    output wire [DATA_WIDTH - 1:0] reg_24_31,
    output wire [DATA_WIDTH - 1:0] reg_29_31,
    output wire [DATA_WIDTH - 1:0] reg_34_31,
    output wire [DATA_WIDTH - 1:0] reg_35_31,
    output wire [DATA_WIDTH - 1:0] reg_16_32,
    output wire [DATA_WIDTH - 1:0] reg_21_32,
    output wire [DATA_WIDTH - 1:0] reg_26_32,
    output wire [DATA_WIDTH - 1:0] reg_27_32,
    output wire [DATA_WIDTH - 1:0] reg_32_32,
    output wire [DATA_WIDTH - 1:0] reg_37_32,
    output wire [DATA_WIDTH - 1:0] reg_14_33,
    output wire [DATA_WIDTH - 1:0] reg_16_33,
    output wire [DATA_WIDTH - 1:0] reg_23_33,
    output wire [DATA_WIDTH - 1:0] reg_30_33,
    output wire [DATA_WIDTH - 1:0] reg_37_33,
    output wire [DATA_WIDTH - 1:0] reg_39_33,
    output wire [DATA_WIDTH - 1:0] reg_12_34,
    output wire [DATA_WIDTH - 1:0] reg_19_34,
    output wire [DATA_WIDTH - 1:0] reg_22_34,
    output wire [DATA_WIDTH - 1:0] reg_26_34,
    output wire [DATA_WIDTH - 1:0] reg_27_34,
    output wire [DATA_WIDTH - 1:0] reg_31_34,
    output wire [DATA_WIDTH - 1:0] reg_34_34,
    output wire [DATA_WIDTH - 1:0] reg_41_34,
    output wire [DATA_WIDTH - 1:0] reg_10_35,
    output wire [DATA_WIDTH - 1:0] reg_13_35,
    output wire [DATA_WIDTH - 1:0] reg_22_35,
    output wire [DATA_WIDTH - 1:0] reg_31_35,
    output wire [DATA_WIDTH - 1:0] reg_40_35,
    output wire [DATA_WIDTH - 1:0] reg_43_35,
    output wire [DATA_WIDTH - 1:0] reg_17_36,
    output wire [DATA_WIDTH - 1:0] reg_26_36,
    output wire [DATA_WIDTH - 1:0] reg_27_36,
    output wire [DATA_WIDTH - 1:0] reg_36_36,
    output wire [DATA_WIDTH - 1:0] reg_10_37,
    output wire [DATA_WIDTH - 1:0] reg_20_37,
    output wire [DATA_WIDTH - 1:0] reg_21_37,
    output wire [DATA_WIDTH - 1:0] reg_32_37,
    output wire [DATA_WIDTH - 1:0] reg_33_37,
    output wire [DATA_WIDTH - 1:0] reg_43_37,
    output wire [DATA_WIDTH - 1:0] reg_15_38,
    output wire [DATA_WIDTH - 1:0] reg_26_38,
    output wire [DATA_WIDTH - 1:0] reg_27_38,
    output wire [DATA_WIDTH - 1:0] reg_38_38,
    output wire [DATA_WIDTH - 1:0] reg_07_39,
    output wire [DATA_WIDTH - 1:0] reg_20_39,
    output wire [DATA_WIDTH - 1:0] reg_33_39,
    output wire [DATA_WIDTH - 1:0] reg_46_39,
    output wire [DATA_WIDTH - 1:0] reg_13_40,
    output wire [DATA_WIDTH - 1:0] reg_18_40,
    output wire [DATA_WIDTH - 1:0] reg_26_40,
    output wire [DATA_WIDTH - 1:0] reg_27_40,
    output wire [DATA_WIDTH - 1:0] reg_35_40,
    output wire [DATA_WIDTH - 1:0] reg_40_40,
    output wire [DATA_WIDTH - 1:0] reg_04_41,
    output wire [DATA_WIDTH - 1:0] reg_19_41,
    output wire [DATA_WIDTH - 1:0] reg_34_41,
    output wire [DATA_WIDTH - 1:0] reg_49_41,
    output wire [DATA_WIDTH - 1:0] reg_11_42,
    output wire [DATA_WIDTH - 1:0] reg_26_42,
    output wire [DATA_WIDTH - 1:0] reg_27_42,
    output wire [DATA_WIDTH - 1:0] reg_42_42,
    output wire [DATA_WIDTH - 1:0] reg_01_43,
    output wire [DATA_WIDTH - 1:0] reg_16_43,
    output wire [DATA_WIDTH - 1:0] reg_18_43,
    output wire [DATA_WIDTH - 1:0] reg_35_43,
    output wire [DATA_WIDTH - 1:0] reg_37_43,
    output wire [DATA_WIDTH - 1:0] reg_52_43,
    output wire [DATA_WIDTH - 1:0] reg_09_44,
    output wire [DATA_WIDTH - 1:0] reg_26_44,
    output wire [DATA_WIDTH - 1:0] reg_27_44,
    output wire [DATA_WIDTH - 1:0] reg_44_44,
    output wire [DATA_WIDTH - 1:0] reg_14_46,
    output wire [DATA_WIDTH - 1:0] reg_39_46,
    output wire [DATA_WIDTH - 1:0] reg_12_49,
    output wire [DATA_WIDTH - 1:0] reg_41_49,
    output wire [DATA_WIDTH - 1:0] reg_10_52,
    output wire [DATA_WIDTH - 1:0] reg_43_52

);

wire [DATA_WIDTH - 1:0] o_d_rowBuf[REGSNUM - 1:1];
wire [DATA_WIDTH - 1:0] o_d_reg[REGSNUM - 1:1][REGSNUM:1];
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH)) rowBuf1
        (
                .din        (din),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[1]),
                .reg01        (o_d_reg[1][1]),
                .reg02        (o_d_reg[1][2]),
                .reg03        (o_d_reg[1][3]),
                .reg04        (o_d_reg[1][4]),
                .reg05        (o_d_reg[1][5]),
                .reg06        (o_d_reg[1][6]),
                .reg07        (o_d_reg[1][7]),
                .reg08        (o_d_reg[1][8]),
                .reg09        (o_d_reg[1][9]),
                .reg10        (o_d_reg[1][10]),
                .reg11        (o_d_reg[1][11]),
                .reg12        (o_d_reg[1][12]),
                .reg13        (o_d_reg[1][13]),
                .reg14        (o_d_reg[1][14]),
                .reg15        (o_d_reg[1][15]),
                .reg16        (o_d_reg[1][16]),
                .reg17        (o_d_reg[1][17]),
                .reg18        (o_d_reg[1][18]),
                .reg19        (o_d_reg[1][19]),
                .reg20        (o_d_reg[1][20]),
                .reg21        (o_d_reg[1][21]),
                .reg22        (o_d_reg[1][22]),
                .reg23        (o_d_reg[1][23]),
                .reg24        (o_d_reg[1][24]),
                .reg25        (o_d_reg[1][25]),
                .reg26        (o_d_reg[1][26]),
                .reg27        (o_d_reg[1][27]),
                .reg28        (o_d_reg[1][28]),
                .reg29        (o_d_reg[1][29]),
                .reg30        (o_d_reg[1][30]),
                .reg31        (o_d_reg[1][31]),
                .reg32        (o_d_reg[1][32]),
                .reg33        (o_d_reg[1][33]),
                .reg34        (o_d_reg[1][34]),
                .reg35        (o_d_reg[1][35]),
                .reg36        (o_d_reg[1][36]),
                .reg37        (o_d_reg[1][37]),
                .reg38        (o_d_reg[1][38]),
                .reg39        (o_d_reg[1][39]),
                .reg40        (o_d_reg[1][40]),
                .reg41        (o_d_reg[1][41]),
                .reg42        (o_d_reg[1][42]),
                .reg43        (o_d_reg[1][43]),
                .reg44        (o_d_reg[1][44]),
                .reg45        (o_d_reg[1][45]),
                .reg46        (o_d_reg[1][46]),
                .reg47        (o_d_reg[1][47]),
                .reg48        (o_d_reg[1][48]),
                .reg49        (o_d_reg[1][49]),
                .reg50        (o_d_reg[1][50]),
                .reg51        (o_d_reg[1][51]),
                .reg52        (o_d_reg[1][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf2
        (
                .din        (o_d_rowBuf[1]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[2]),
                .reg01        (o_d_reg[2][1]),
                .reg02        (o_d_reg[2][2]),
                .reg03        (o_d_reg[2][3]),
                .reg04        (o_d_reg[2][4]),
                .reg05        (o_d_reg[2][5]),
                .reg06        (o_d_reg[2][6]),
                .reg07        (o_d_reg[2][7]),
                .reg08        (o_d_reg[2][8]),
                .reg09        (o_d_reg[2][9]),
                .reg10        (o_d_reg[2][10]),
                .reg11        (o_d_reg[2][11]),
                .reg12        (o_d_reg[2][12]),
                .reg13        (o_d_reg[2][13]),
                .reg14        (o_d_reg[2][14]),
                .reg15        (o_d_reg[2][15]),
                .reg16        (o_d_reg[2][16]),
                .reg17        (o_d_reg[2][17]),
                .reg18        (o_d_reg[2][18]),
                .reg19        (o_d_reg[2][19]),
                .reg20        (o_d_reg[2][20]),
                .reg21        (o_d_reg[2][21]),
                .reg22        (o_d_reg[2][22]),
                .reg23        (o_d_reg[2][23]),
                .reg24        (o_d_reg[2][24]),
                .reg25        (o_d_reg[2][25]),
                .reg26        (o_d_reg[2][26]),
                .reg27        (o_d_reg[2][27]),
                .reg28        (o_d_reg[2][28]),
                .reg29        (o_d_reg[2][29]),
                .reg30        (o_d_reg[2][30]),
                .reg31        (o_d_reg[2][31]),
                .reg32        (o_d_reg[2][32]),
                .reg33        (o_d_reg[2][33]),
                .reg34        (o_d_reg[2][34]),
                .reg35        (o_d_reg[2][35]),
                .reg36        (o_d_reg[2][36]),
                .reg37        (o_d_reg[2][37]),
                .reg38        (o_d_reg[2][38]),
                .reg39        (o_d_reg[2][39]),
                .reg40        (o_d_reg[2][40]),
                .reg41        (o_d_reg[2][41]),
                .reg42        (o_d_reg[2][42]),
                .reg43        (o_d_reg[2][43]),
                .reg44        (o_d_reg[2][44]),
                .reg45        (o_d_reg[2][45]),
                .reg46        (o_d_reg[2][46]),
                .reg47        (o_d_reg[2][47]),
                .reg48        (o_d_reg[2][48]),
                .reg49        (o_d_reg[2][49]),
                .reg50        (o_d_reg[2][50]),
                .reg51        (o_d_reg[2][51]),
                .reg52        (o_d_reg[2][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf3
        (
                .din        (o_d_rowBuf[2]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[3]),
                .reg01        (o_d_reg[3][1]),
                .reg02        (o_d_reg[3][2]),
                .reg03        (o_d_reg[3][3]),
                .reg04        (o_d_reg[3][4]),
                .reg05        (o_d_reg[3][5]),
                .reg06        (o_d_reg[3][6]),
                .reg07        (o_d_reg[3][7]),
                .reg08        (o_d_reg[3][8]),
                .reg09        (o_d_reg[3][9]),
                .reg10        (o_d_reg[3][10]),
                .reg11        (o_d_reg[3][11]),
                .reg12        (o_d_reg[3][12]),
                .reg13        (o_d_reg[3][13]),
                .reg14        (o_d_reg[3][14]),
                .reg15        (o_d_reg[3][15]),
                .reg16        (o_d_reg[3][16]),
                .reg17        (o_d_reg[3][17]),
                .reg18        (o_d_reg[3][18]),
                .reg19        (o_d_reg[3][19]),
                .reg20        (o_d_reg[3][20]),
                .reg21        (o_d_reg[3][21]),
                .reg22        (o_d_reg[3][22]),
                .reg23        (o_d_reg[3][23]),
                .reg24        (o_d_reg[3][24]),
                .reg25        (o_d_reg[3][25]),
                .reg26        (o_d_reg[3][26]),
                .reg27        (o_d_reg[3][27]),
                .reg28        (o_d_reg[3][28]),
                .reg29        (o_d_reg[3][29]),
                .reg30        (o_d_reg[3][30]),
                .reg31        (o_d_reg[3][31]),
                .reg32        (o_d_reg[3][32]),
                .reg33        (o_d_reg[3][33]),
                .reg34        (o_d_reg[3][34]),
                .reg35        (o_d_reg[3][35]),
                .reg36        (o_d_reg[3][36]),
                .reg37        (o_d_reg[3][37]),
                .reg38        (o_d_reg[3][38]),
                .reg39        (o_d_reg[3][39]),
                .reg40        (o_d_reg[3][40]),
                .reg41        (o_d_reg[3][41]),
                .reg42        (o_d_reg[3][42]),
                .reg43        (o_d_reg[3][43]),
                .reg44        (o_d_reg[3][44]),
                .reg45        (o_d_reg[3][45]),
                .reg46        (o_d_reg[3][46]),
                .reg47        (o_d_reg[3][47]),
                .reg48        (o_d_reg[3][48]),
                .reg49        (o_d_reg[3][49]),
                .reg50        (o_d_reg[3][50]),
                .reg51        (o_d_reg[3][51]),
                .reg52        (o_d_reg[3][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf4
        (
                .din        (o_d_rowBuf[3]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[4]),
                .reg01        (o_d_reg[4][1]),
                .reg02        (o_d_reg[4][2]),
                .reg03        (o_d_reg[4][3]),
                .reg04        (o_d_reg[4][4]),
                .reg05        (o_d_reg[4][5]),
                .reg06        (o_d_reg[4][6]),
                .reg07        (o_d_reg[4][7]),
                .reg08        (o_d_reg[4][8]),
                .reg09        (o_d_reg[4][9]),
                .reg10        (o_d_reg[4][10]),
                .reg11        (o_d_reg[4][11]),
                .reg12        (o_d_reg[4][12]),
                .reg13        (o_d_reg[4][13]),
                .reg14        (o_d_reg[4][14]),
                .reg15        (o_d_reg[4][15]),
                .reg16        (o_d_reg[4][16]),
                .reg17        (o_d_reg[4][17]),
                .reg18        (o_d_reg[4][18]),
                .reg19        (o_d_reg[4][19]),
                .reg20        (o_d_reg[4][20]),
                .reg21        (o_d_reg[4][21]),
                .reg22        (o_d_reg[4][22]),
                .reg23        (o_d_reg[4][23]),
                .reg24        (o_d_reg[4][24]),
                .reg25        (o_d_reg[4][25]),
                .reg26        (o_d_reg[4][26]),
                .reg27        (o_d_reg[4][27]),
                .reg28        (o_d_reg[4][28]),
                .reg29        (o_d_reg[4][29]),
                .reg30        (o_d_reg[4][30]),
                .reg31        (o_d_reg[4][31]),
                .reg32        (o_d_reg[4][32]),
                .reg33        (o_d_reg[4][33]),
                .reg34        (o_d_reg[4][34]),
                .reg35        (o_d_reg[4][35]),
                .reg36        (o_d_reg[4][36]),
                .reg37        (o_d_reg[4][37]),
                .reg38        (o_d_reg[4][38]),
                .reg39        (o_d_reg[4][39]),
                .reg40        (o_d_reg[4][40]),
                .reg41        (o_d_reg[4][41]),
                .reg42        (o_d_reg[4][42]),
                .reg43        (o_d_reg[4][43]),
                .reg44        (o_d_reg[4][44]),
                .reg45        (o_d_reg[4][45]),
                .reg46        (o_d_reg[4][46]),
                .reg47        (o_d_reg[4][47]),
                .reg48        (o_d_reg[4][48]),
                .reg49        (o_d_reg[4][49]),
                .reg50        (o_d_reg[4][50]),
                .reg51        (o_d_reg[4][51]),
                .reg52        (o_d_reg[4][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf5
        (
                .din        (o_d_rowBuf[4]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[5]),
                .reg01        (o_d_reg[5][1]),
                .reg02        (o_d_reg[5][2]),
                .reg03        (o_d_reg[5][3]),
                .reg04        (o_d_reg[5][4]),
                .reg05        (o_d_reg[5][5]),
                .reg06        (o_d_reg[5][6]),
                .reg07        (o_d_reg[5][7]),
                .reg08        (o_d_reg[5][8]),
                .reg09        (o_d_reg[5][9]),
                .reg10        (o_d_reg[5][10]),
                .reg11        (o_d_reg[5][11]),
                .reg12        (o_d_reg[5][12]),
                .reg13        (o_d_reg[5][13]),
                .reg14        (o_d_reg[5][14]),
                .reg15        (o_d_reg[5][15]),
                .reg16        (o_d_reg[5][16]),
                .reg17        (o_d_reg[5][17]),
                .reg18        (o_d_reg[5][18]),
                .reg19        (o_d_reg[5][19]),
                .reg20        (o_d_reg[5][20]),
                .reg21        (o_d_reg[5][21]),
                .reg22        (o_d_reg[5][22]),
                .reg23        (o_d_reg[5][23]),
                .reg24        (o_d_reg[5][24]),
                .reg25        (o_d_reg[5][25]),
                .reg26        (o_d_reg[5][26]),
                .reg27        (o_d_reg[5][27]),
                .reg28        (o_d_reg[5][28]),
                .reg29        (o_d_reg[5][29]),
                .reg30        (o_d_reg[5][30]),
                .reg31        (o_d_reg[5][31]),
                .reg32        (o_d_reg[5][32]),
                .reg33        (o_d_reg[5][33]),
                .reg34        (o_d_reg[5][34]),
                .reg35        (o_d_reg[5][35]),
                .reg36        (o_d_reg[5][36]),
                .reg37        (o_d_reg[5][37]),
                .reg38        (o_d_reg[5][38]),
                .reg39        (o_d_reg[5][39]),
                .reg40        (o_d_reg[5][40]),
                .reg41        (o_d_reg[5][41]),
                .reg42        (o_d_reg[5][42]),
                .reg43        (o_d_reg[5][43]),
                .reg44        (o_d_reg[5][44]),
                .reg45        (o_d_reg[5][45]),
                .reg46        (o_d_reg[5][46]),
                .reg47        (o_d_reg[5][47]),
                .reg48        (o_d_reg[5][48]),
                .reg49        (o_d_reg[5][49]),
                .reg50        (o_d_reg[5][50]),
                .reg51        (o_d_reg[5][51]),
                .reg52        (o_d_reg[5][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf6
        (
                .din        (o_d_rowBuf[5]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[6]),
                .reg01        (o_d_reg[6][1]),
                .reg02        (o_d_reg[6][2]),
                .reg03        (o_d_reg[6][3]),
                .reg04        (o_d_reg[6][4]),
                .reg05        (o_d_reg[6][5]),
                .reg06        (o_d_reg[6][6]),
                .reg07        (o_d_reg[6][7]),
                .reg08        (o_d_reg[6][8]),
                .reg09        (o_d_reg[6][9]),
                .reg10        (o_d_reg[6][10]),
                .reg11        (o_d_reg[6][11]),
                .reg12        (o_d_reg[6][12]),
                .reg13        (o_d_reg[6][13]),
                .reg14        (o_d_reg[6][14]),
                .reg15        (o_d_reg[6][15]),
                .reg16        (o_d_reg[6][16]),
                .reg17        (o_d_reg[6][17]),
                .reg18        (o_d_reg[6][18]),
                .reg19        (o_d_reg[6][19]),
                .reg20        (o_d_reg[6][20]),
                .reg21        (o_d_reg[6][21]),
                .reg22        (o_d_reg[6][22]),
                .reg23        (o_d_reg[6][23]),
                .reg24        (o_d_reg[6][24]),
                .reg25        (o_d_reg[6][25]),
                .reg26        (o_d_reg[6][26]),
                .reg27        (o_d_reg[6][27]),
                .reg28        (o_d_reg[6][28]),
                .reg29        (o_d_reg[6][29]),
                .reg30        (o_d_reg[6][30]),
                .reg31        (o_d_reg[6][31]),
                .reg32        (o_d_reg[6][32]),
                .reg33        (o_d_reg[6][33]),
                .reg34        (o_d_reg[6][34]),
                .reg35        (o_d_reg[6][35]),
                .reg36        (o_d_reg[6][36]),
                .reg37        (o_d_reg[6][37]),
                .reg38        (o_d_reg[6][38]),
                .reg39        (o_d_reg[6][39]),
                .reg40        (o_d_reg[6][40]),
                .reg41        (o_d_reg[6][41]),
                .reg42        (o_d_reg[6][42]),
                .reg43        (o_d_reg[6][43]),
                .reg44        (o_d_reg[6][44]),
                .reg45        (o_d_reg[6][45]),
                .reg46        (o_d_reg[6][46]),
                .reg47        (o_d_reg[6][47]),
                .reg48        (o_d_reg[6][48]),
                .reg49        (o_d_reg[6][49]),
                .reg50        (o_d_reg[6][50]),
                .reg51        (o_d_reg[6][51]),
                .reg52        (o_d_reg[6][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf7
        (
                .din        (o_d_rowBuf[6]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[7]),
                .reg01        (o_d_reg[7][1]),
                .reg02        (o_d_reg[7][2]),
                .reg03        (o_d_reg[7][3]),
                .reg04        (o_d_reg[7][4]),
                .reg05        (o_d_reg[7][5]),
                .reg06        (o_d_reg[7][6]),
                .reg07        (o_d_reg[7][7]),
                .reg08        (o_d_reg[7][8]),
                .reg09        (o_d_reg[7][9]),
                .reg10        (o_d_reg[7][10]),
                .reg11        (o_d_reg[7][11]),
                .reg12        (o_d_reg[7][12]),
                .reg13        (o_d_reg[7][13]),
                .reg14        (o_d_reg[7][14]),
                .reg15        (o_d_reg[7][15]),
                .reg16        (o_d_reg[7][16]),
                .reg17        (o_d_reg[7][17]),
                .reg18        (o_d_reg[7][18]),
                .reg19        (o_d_reg[7][19]),
                .reg20        (o_d_reg[7][20]),
                .reg21        (o_d_reg[7][21]),
                .reg22        (o_d_reg[7][22]),
                .reg23        (o_d_reg[7][23]),
                .reg24        (o_d_reg[7][24]),
                .reg25        (o_d_reg[7][25]),
                .reg26        (o_d_reg[7][26]),
                .reg27        (o_d_reg[7][27]),
                .reg28        (o_d_reg[7][28]),
                .reg29        (o_d_reg[7][29]),
                .reg30        (o_d_reg[7][30]),
                .reg31        (o_d_reg[7][31]),
                .reg32        (o_d_reg[7][32]),
                .reg33        (o_d_reg[7][33]),
                .reg34        (o_d_reg[7][34]),
                .reg35        (o_d_reg[7][35]),
                .reg36        (o_d_reg[7][36]),
                .reg37        (o_d_reg[7][37]),
                .reg38        (o_d_reg[7][38]),
                .reg39        (o_d_reg[7][39]),
                .reg40        (o_d_reg[7][40]),
                .reg41        (o_d_reg[7][41]),
                .reg42        (o_d_reg[7][42]),
                .reg43        (o_d_reg[7][43]),
                .reg44        (o_d_reg[7][44]),
                .reg45        (o_d_reg[7][45]),
                .reg46        (o_d_reg[7][46]),
                .reg47        (o_d_reg[7][47]),
                .reg48        (o_d_reg[7][48]),
                .reg49        (o_d_reg[7][49]),
                .reg50        (o_d_reg[7][50]),
                .reg51        (o_d_reg[7][51]),
                .reg52        (o_d_reg[7][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf8
        (
                .din        (o_d_rowBuf[7]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[8]),
                .reg01        (o_d_reg[8][1]),
                .reg02        (o_d_reg[8][2]),
                .reg03        (o_d_reg[8][3]),
                .reg04        (o_d_reg[8][4]),
                .reg05        (o_d_reg[8][5]),
                .reg06        (o_d_reg[8][6]),
                .reg07        (o_d_reg[8][7]),
                .reg08        (o_d_reg[8][8]),
                .reg09        (o_d_reg[8][9]),
                .reg10        (o_d_reg[8][10]),
                .reg11        (o_d_reg[8][11]),
                .reg12        (o_d_reg[8][12]),
                .reg13        (o_d_reg[8][13]),
                .reg14        (o_d_reg[8][14]),
                .reg15        (o_d_reg[8][15]),
                .reg16        (o_d_reg[8][16]),
                .reg17        (o_d_reg[8][17]),
                .reg18        (o_d_reg[8][18]),
                .reg19        (o_d_reg[8][19]),
                .reg20        (o_d_reg[8][20]),
                .reg21        (o_d_reg[8][21]),
                .reg22        (o_d_reg[8][22]),
                .reg23        (o_d_reg[8][23]),
                .reg24        (o_d_reg[8][24]),
                .reg25        (o_d_reg[8][25]),
                .reg26        (o_d_reg[8][26]),
                .reg27        (o_d_reg[8][27]),
                .reg28        (o_d_reg[8][28]),
                .reg29        (o_d_reg[8][29]),
                .reg30        (o_d_reg[8][30]),
                .reg31        (o_d_reg[8][31]),
                .reg32        (o_d_reg[8][32]),
                .reg33        (o_d_reg[8][33]),
                .reg34        (o_d_reg[8][34]),
                .reg35        (o_d_reg[8][35]),
                .reg36        (o_d_reg[8][36]),
                .reg37        (o_d_reg[8][37]),
                .reg38        (o_d_reg[8][38]),
                .reg39        (o_d_reg[8][39]),
                .reg40        (o_d_reg[8][40]),
                .reg41        (o_d_reg[8][41]),
                .reg42        (o_d_reg[8][42]),
                .reg43        (o_d_reg[8][43]),
                .reg44        (o_d_reg[8][44]),
                .reg45        (o_d_reg[8][45]),
                .reg46        (o_d_reg[8][46]),
                .reg47        (o_d_reg[8][47]),
                .reg48        (o_d_reg[8][48]),
                .reg49        (o_d_reg[8][49]),
                .reg50        (o_d_reg[8][50]),
                .reg51        (o_d_reg[8][51]),
                .reg52        (o_d_reg[8][52])
        );

        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf9
        (
                .din        (o_d_rowBuf[8]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[9]),
                .reg01        (o_d_reg[9][1]),
                .reg02        (o_d_reg[9][2]),
                .reg03        (o_d_reg[9][3]),
                .reg04        (o_d_reg[9][4]),
                .reg05        (o_d_reg[9][5]),
                .reg06        (o_d_reg[9][6]),
                .reg07        (o_d_reg[9][7]),
                .reg08        (o_d_reg[9][8]),
                .reg09        (o_d_reg[9][9]),
                .reg10        (o_d_reg[9][10]),
                .reg11        (o_d_reg[9][11]),
                .reg12        (o_d_reg[9][12]),
                .reg13        (o_d_reg[9][13]),
                .reg14        (o_d_reg[9][14]),
                .reg15        (o_d_reg[9][15]),
                .reg16        (o_d_reg[9][16]),
                .reg17        (o_d_reg[9][17]),
                .reg18        (o_d_reg[9][18]),
                .reg19        (o_d_reg[9][19]),
                .reg20        (o_d_reg[9][20]),
                .reg21        (o_d_reg[9][21]),
                .reg22        (o_d_reg[9][22]),
                .reg23        (o_d_reg[9][23]),
                .reg24        (o_d_reg[9][24]),
                .reg25        (o_d_reg[9][25]),
                .reg26        (o_d_reg[9][26]),
                .reg27        (o_d_reg[9][27]),
                .reg28        (o_d_reg[9][28]),
                .reg29        (o_d_reg[9][29]),
                .reg30        (o_d_reg[9][30]),
                .reg31        (o_d_reg[9][31]),
                .reg32        (o_d_reg[9][32]),
                .reg33        (o_d_reg[9][33]),
                .reg34        (o_d_reg[9][34]),
                .reg35        (o_d_reg[9][35]),
                .reg36        (o_d_reg[9][36]),
                .reg37        (o_d_reg[9][37]),
                .reg38        (o_d_reg[9][38]),
                .reg39        (o_d_reg[9][39]),
                .reg40        (o_d_reg[9][40]),
                .reg41        (o_d_reg[9][41]),
                .reg42        (o_d_reg[9][42]),
                .reg43        (o_d_reg[9][43]),
                .reg44        (o_d_reg[9][44]),
                .reg45        (o_d_reg[9][45]),
                .reg46        (o_d_reg[9][46]),
                .reg47        (o_d_reg[9][47]),
                .reg48        (o_d_reg[9][48]),
                .reg49        (o_d_reg[9][49]),
                .reg50        (o_d_reg[9][50]),
                .reg51        (o_d_reg[9][51]),
                .reg52        (o_d_reg[9][52])
        );		
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf10
        (
                .din        (o_d_rowBuf[9]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[10]),
                .reg01        (o_d_reg[10][1]),
                .reg02        (o_d_reg[10][2]),
                .reg03        (o_d_reg[10][3]),
                .reg04        (o_d_reg[10][4]),
                .reg05        (o_d_reg[10][5]),
                .reg06        (o_d_reg[10][6]),
                .reg07        (o_d_reg[10][7]),
                .reg08        (o_d_reg[10][8]),
                .reg09        (o_d_reg[10][9]),
                .reg10        (o_d_reg[10][10]),
                .reg11        (o_d_reg[10][11]),
                .reg12        (o_d_reg[10][12]),
                .reg13        (o_d_reg[10][13]),
                .reg14        (o_d_reg[10][14]),
                .reg15        (o_d_reg[10][15]),
                .reg16        (o_d_reg[10][16]),
                .reg17        (o_d_reg[10][17]),
                .reg18        (o_d_reg[10][18]),
                .reg19        (o_d_reg[10][19]),
                .reg20        (o_d_reg[10][20]),
                .reg21        (o_d_reg[10][21]),
                .reg22        (o_d_reg[10][22]),
                .reg23        (o_d_reg[10][23]),
                .reg24        (o_d_reg[10][24]),
                .reg25        (o_d_reg[10][25]),
                .reg26        (o_d_reg[10][26]),
                .reg27        (o_d_reg[10][27]),
                .reg28        (o_d_reg[10][28]),
                .reg29        (o_d_reg[10][29]),
                .reg30        (o_d_reg[10][30]),
                .reg31        (o_d_reg[10][31]),
                .reg32        (o_d_reg[10][32]),
                .reg33        (o_d_reg[10][33]),
                .reg34        (o_d_reg[10][34]),
                .reg35        (o_d_reg[10][35]),
                .reg36        (o_d_reg[10][36]),
                .reg37        (o_d_reg[10][37]),
                .reg38        (o_d_reg[10][38]),
                .reg39        (o_d_reg[10][39]),
                .reg40        (o_d_reg[10][40]),
                .reg41        (o_d_reg[10][41]),
                .reg42        (o_d_reg[10][42]),
                .reg43        (o_d_reg[10][43]),
                .reg44        (o_d_reg[10][44]),
                .reg45        (o_d_reg[10][45]),
                .reg46        (o_d_reg[10][46]),
                .reg47        (o_d_reg[10][47]),
                .reg48        (o_d_reg[10][48]),
                .reg49        (o_d_reg[10][49]),
                .reg50        (o_d_reg[10][50]),
                .reg51        (o_d_reg[10][51]),
                .reg52        (o_d_reg[10][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf11
        (
                .din        (o_d_rowBuf[10]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[11]),
                .reg01        (o_d_reg[11][1]),
                .reg02        (o_d_reg[11][2]),
                .reg03        (o_d_reg[11][3]),
                .reg04        (o_d_reg[11][4]),
                .reg05        (o_d_reg[11][5]),
                .reg06        (o_d_reg[11][6]),
                .reg07        (o_d_reg[11][7]),
                .reg08        (o_d_reg[11][8]),
                .reg09        (o_d_reg[11][9]),
                .reg10        (o_d_reg[11][10]),
                .reg11        (o_d_reg[11][11]),
                .reg12        (o_d_reg[11][12]),
                .reg13        (o_d_reg[11][13]),
                .reg14        (o_d_reg[11][14]),
                .reg15        (o_d_reg[11][15]),
                .reg16        (o_d_reg[11][16]),
                .reg17        (o_d_reg[11][17]),
                .reg18        (o_d_reg[11][18]),
                .reg19        (o_d_reg[11][19]),
                .reg20        (o_d_reg[11][20]),
                .reg21        (o_d_reg[11][21]),
                .reg22        (o_d_reg[11][22]),
                .reg23        (o_d_reg[11][23]),
                .reg24        (o_d_reg[11][24]),
                .reg25        (o_d_reg[11][25]),
                .reg26        (o_d_reg[11][26]),
                .reg27        (o_d_reg[11][27]),
                .reg28        (o_d_reg[11][28]),
                .reg29        (o_d_reg[11][29]),
                .reg30        (o_d_reg[11][30]),
                .reg31        (o_d_reg[11][31]),
                .reg32        (o_d_reg[11][32]),
                .reg33        (o_d_reg[11][33]),
                .reg34        (o_d_reg[11][34]),
                .reg35        (o_d_reg[11][35]),
                .reg36        (o_d_reg[11][36]),
                .reg37        (o_d_reg[11][37]),
                .reg38        (o_d_reg[11][38]),
                .reg39        (o_d_reg[11][39]),
                .reg40        (o_d_reg[11][40]),
                .reg41        (o_d_reg[11][41]),
                .reg42        (o_d_reg[11][42]),
                .reg43        (o_d_reg[11][43]),
                .reg44        (o_d_reg[11][44]),
                .reg45        (o_d_reg[11][45]),
                .reg46        (o_d_reg[11][46]),
                .reg47        (o_d_reg[11][47]),
                .reg48        (o_d_reg[11][48]),
                .reg49        (o_d_reg[11][49]),
                .reg50        (o_d_reg[11][50]),
                .reg51        (o_d_reg[11][51]),
                .reg52        (o_d_reg[11][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf12
        (
                .din        (o_d_rowBuf[11]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[12]),
                .reg01        (o_d_reg[12][1]),
                .reg02        (o_d_reg[12][2]),
                .reg03        (o_d_reg[12][3]),
                .reg04        (o_d_reg[12][4]),
                .reg05        (o_d_reg[12][5]),
                .reg06        (o_d_reg[12][6]),
                .reg07        (o_d_reg[12][7]),
                .reg08        (o_d_reg[12][8]),
                .reg09        (o_d_reg[12][9]),
                .reg10        (o_d_reg[12][10]),
                .reg11        (o_d_reg[12][11]),
                .reg12        (o_d_reg[12][12]),
                .reg13        (o_d_reg[12][13]),
                .reg14        (o_d_reg[12][14]),
                .reg15        (o_d_reg[12][15]),
                .reg16        (o_d_reg[12][16]),
                .reg17        (o_d_reg[12][17]),
                .reg18        (o_d_reg[12][18]),
                .reg19        (o_d_reg[12][19]),
                .reg20        (o_d_reg[12][20]),
                .reg21        (o_d_reg[12][21]),
                .reg22        (o_d_reg[12][22]),
                .reg23        (o_d_reg[12][23]),
                .reg24        (o_d_reg[12][24]),
                .reg25        (o_d_reg[12][25]),
                .reg26        (o_d_reg[12][26]),
                .reg27        (o_d_reg[12][27]),
                .reg28        (o_d_reg[12][28]),
                .reg29        (o_d_reg[12][29]),
                .reg30        (o_d_reg[12][30]),
                .reg31        (o_d_reg[12][31]),
                .reg32        (o_d_reg[12][32]),
                .reg33        (o_d_reg[12][33]),
                .reg34        (o_d_reg[12][34]),
                .reg35        (o_d_reg[12][35]),
                .reg36        (o_d_reg[12][36]),
                .reg37        (o_d_reg[12][37]),
                .reg38        (o_d_reg[12][38]),
                .reg39        (o_d_reg[12][39]),
                .reg40        (o_d_reg[12][40]),
                .reg41        (o_d_reg[12][41]),
                .reg42        (o_d_reg[12][42]),
                .reg43        (o_d_reg[12][43]),
                .reg44        (o_d_reg[12][44]),
                .reg45        (o_d_reg[12][45]),
                .reg46        (o_d_reg[12][46]),
                .reg47        (o_d_reg[12][47]),
                .reg48        (o_d_reg[12][48]),
                .reg49        (o_d_reg[12][49]),
                .reg50        (o_d_reg[12][50]),
                .reg51        (o_d_reg[12][51]),
                .reg52        (o_d_reg[12][52])
        );	
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf13
        (
                .din        (o_d_rowBuf[12]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[13]),
                .reg01        (o_d_reg[13][1]),
                .reg02        (o_d_reg[13][2]),
                .reg03        (o_d_reg[13][3]),
                .reg04        (o_d_reg[13][4]),
                .reg05        (o_d_reg[13][5]),
                .reg06        (o_d_reg[13][6]),
                .reg07        (o_d_reg[13][7]),
                .reg08        (o_d_reg[13][8]),
                .reg09        (o_d_reg[13][9]),
                .reg10        (o_d_reg[13][10]),
                .reg11        (o_d_reg[13][11]),
                .reg12        (o_d_reg[13][12]),
                .reg13        (o_d_reg[13][13]),
                .reg14        (o_d_reg[13][14]),
                .reg15        (o_d_reg[13][15]),
                .reg16        (o_d_reg[13][16]),
                .reg17        (o_d_reg[13][17]),
                .reg18        (o_d_reg[13][18]),
                .reg19        (o_d_reg[13][19]),
                .reg20        (o_d_reg[13][20]),
                .reg21        (o_d_reg[13][21]),
                .reg22        (o_d_reg[13][22]),
                .reg23        (o_d_reg[13][23]),
                .reg24        (o_d_reg[13][24]),
                .reg25        (o_d_reg[13][25]),
                .reg26        (o_d_reg[13][26]),
                .reg27        (o_d_reg[13][27]),
                .reg28        (o_d_reg[13][28]),
                .reg29        (o_d_reg[13][29]),
                .reg30        (o_d_reg[13][30]),
                .reg31        (o_d_reg[13][31]),
                .reg32        (o_d_reg[13][32]),
                .reg33        (o_d_reg[13][33]),
                .reg34        (o_d_reg[13][34]),
                .reg35        (o_d_reg[13][35]),
                .reg36        (o_d_reg[13][36]),
                .reg37        (o_d_reg[13][37]),
                .reg38        (o_d_reg[13][38]),
                .reg39        (o_d_reg[13][39]),
                .reg40        (o_d_reg[13][40]),
                .reg41        (o_d_reg[13][41]),
                .reg42        (o_d_reg[13][42]),
                .reg43        (o_d_reg[13][43]),
                .reg44        (o_d_reg[13][44]),
                .reg45        (o_d_reg[13][45]),
                .reg46        (o_d_reg[13][46]),
                .reg47        (o_d_reg[13][47]),
                .reg48        (o_d_reg[13][48]),
                .reg49        (o_d_reg[13][49]),
                .reg50        (o_d_reg[13][50]),
                .reg51        (o_d_reg[13][51]),
                .reg52        (o_d_reg[13][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf14
        (
                .din        (o_d_rowBuf[13]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[14]),
                .reg01        (o_d_reg[14][1]),
                .reg02        (o_d_reg[14][2]),
                .reg03        (o_d_reg[14][3]),
                .reg04        (o_d_reg[14][4]),
                .reg05        (o_d_reg[14][5]),
                .reg06        (o_d_reg[14][6]),
                .reg07        (o_d_reg[14][7]),
                .reg08        (o_d_reg[14][8]),
                .reg09        (o_d_reg[14][9]),
                .reg10        (o_d_reg[14][10]),
                .reg11        (o_d_reg[14][11]),
                .reg12        (o_d_reg[14][12]),
                .reg13        (o_d_reg[14][13]),
                .reg14        (o_d_reg[14][14]),
                .reg15        (o_d_reg[14][15]),
                .reg16        (o_d_reg[14][16]),
                .reg17        (o_d_reg[14][17]),
                .reg18        (o_d_reg[14][18]),
                .reg19        (o_d_reg[14][19]),
                .reg20        (o_d_reg[14][20]),
                .reg21        (o_d_reg[14][21]),
                .reg22        (o_d_reg[14][22]),
                .reg23        (o_d_reg[14][23]),
                .reg24        (o_d_reg[14][24]),
                .reg25        (o_d_reg[14][25]),
                .reg26        (o_d_reg[14][26]),
                .reg27        (o_d_reg[14][27]),
                .reg28        (o_d_reg[14][28]),
                .reg29        (o_d_reg[14][29]),
                .reg30        (o_d_reg[14][30]),
                .reg31        (o_d_reg[14][31]),
                .reg32        (o_d_reg[14][32]),
                .reg33        (o_d_reg[14][33]),
                .reg34        (o_d_reg[14][34]),
                .reg35        (o_d_reg[14][35]),
                .reg36        (o_d_reg[14][36]),
                .reg37        (o_d_reg[14][37]),
                .reg38        (o_d_reg[14][38]),
                .reg39        (o_d_reg[14][39]),
                .reg40        (o_d_reg[14][40]),
                .reg41        (o_d_reg[14][41]),
                .reg42        (o_d_reg[14][42]),
                .reg43        (o_d_reg[14][43]),
                .reg44        (o_d_reg[14][44]),
                .reg45        (o_d_reg[14][45]),
                .reg46        (o_d_reg[14][46]),
                .reg47        (o_d_reg[14][47]),
                .reg48        (o_d_reg[14][48]),
                .reg49        (o_d_reg[14][49]),
                .reg50        (o_d_reg[14][50]),
                .reg51        (o_d_reg[14][51]),
                .reg52        (o_d_reg[14][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf15
        (
                .din        (o_d_rowBuf[14]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[15]),
                .reg01        (o_d_reg[15][1]),
                .reg02        (o_d_reg[15][2]),
                .reg03        (o_d_reg[15][3]),
                .reg04        (o_d_reg[15][4]),
                .reg05        (o_d_reg[15][5]),
                .reg06        (o_d_reg[15][6]),
                .reg07        (o_d_reg[15][7]),
                .reg08        (o_d_reg[15][8]),
                .reg09        (o_d_reg[15][9]),
                .reg10        (o_d_reg[15][10]),
                .reg11        (o_d_reg[15][11]),
                .reg12        (o_d_reg[15][12]),
                .reg13        (o_d_reg[15][13]),
                .reg14        (o_d_reg[15][14]),
                .reg15        (o_d_reg[15][15]),
                .reg16        (o_d_reg[15][16]),
                .reg17        (o_d_reg[15][17]),
                .reg18        (o_d_reg[15][18]),
                .reg19        (o_d_reg[15][19]),
                .reg20        (o_d_reg[15][20]),
                .reg21        (o_d_reg[15][21]),
                .reg22        (o_d_reg[15][22]),
                .reg23        (o_d_reg[15][23]),
                .reg24        (o_d_reg[15][24]),
                .reg25        (o_d_reg[15][25]),
                .reg26        (o_d_reg[15][26]),
                .reg27        (o_d_reg[15][27]),
                .reg28        (o_d_reg[15][28]),
                .reg29        (o_d_reg[15][29]),
                .reg30        (o_d_reg[15][30]),
                .reg31        (o_d_reg[15][31]),
                .reg32        (o_d_reg[15][32]),
                .reg33        (o_d_reg[15][33]),
                .reg34        (o_d_reg[15][34]),
                .reg35        (o_d_reg[15][35]),
                .reg36        (o_d_reg[15][36]),
                .reg37        (o_d_reg[15][37]),
                .reg38        (o_d_reg[15][38]),
                .reg39        (o_d_reg[15][39]),
                .reg40        (o_d_reg[15][40]),
                .reg41        (o_d_reg[15][41]),
                .reg42        (o_d_reg[15][42]),
                .reg43        (o_d_reg[15][43]),
                .reg44        (o_d_reg[15][44]),
                .reg45        (o_d_reg[15][45]),
                .reg46        (o_d_reg[15][46]),
                .reg47        (o_d_reg[15][47]),
                .reg48        (o_d_reg[15][48]),
                .reg49        (o_d_reg[15][49]),
                .reg50        (o_d_reg[15][50]),
                .reg51        (o_d_reg[15][51]),
                .reg52        (o_d_reg[15][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf16
        (
                .din        (o_d_rowBuf[15]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[16]),
                .reg01        (o_d_reg[16][1]),
                .reg02        (o_d_reg[16][2]),
                .reg03        (o_d_reg[16][3]),
                .reg04        (o_d_reg[16][4]),
                .reg05        (o_d_reg[16][5]),
                .reg06        (o_d_reg[16][6]),
                .reg07        (o_d_reg[16][7]),
                .reg08        (o_d_reg[16][8]),
                .reg09        (o_d_reg[16][9]),
                .reg10        (o_d_reg[16][10]),
                .reg11        (o_d_reg[16][11]),
                .reg12        (o_d_reg[16][12]),
                .reg13        (o_d_reg[16][13]),
                .reg14        (o_d_reg[16][14]),
                .reg15        (o_d_reg[16][15]),
                .reg16        (o_d_reg[16][16]),
                .reg17        (o_d_reg[16][17]),
                .reg18        (o_d_reg[16][18]),
                .reg19        (o_d_reg[16][19]),
                .reg20        (o_d_reg[16][20]),
                .reg21        (o_d_reg[16][21]),
                .reg22        (o_d_reg[16][22]),
                .reg23        (o_d_reg[16][23]),
                .reg24        (o_d_reg[16][24]),
                .reg25        (o_d_reg[16][25]),
                .reg26        (o_d_reg[16][26]),
                .reg27        (o_d_reg[16][27]),
                .reg28        (o_d_reg[16][28]),
                .reg29        (o_d_reg[16][29]),
                .reg30        (o_d_reg[16][30]),
                .reg31        (o_d_reg[16][31]),
                .reg32        (o_d_reg[16][32]),
                .reg33        (o_d_reg[16][33]),
                .reg34        (o_d_reg[16][34]),
                .reg35        (o_d_reg[16][35]),
                .reg36        (o_d_reg[16][36]),
                .reg37        (o_d_reg[16][37]),
                .reg38        (o_d_reg[16][38]),
                .reg39        (o_d_reg[16][39]),
                .reg40        (o_d_reg[16][40]),
                .reg41        (o_d_reg[16][41]),
                .reg42        (o_d_reg[16][42]),
                .reg43        (o_d_reg[16][43]),
                .reg44        (o_d_reg[16][44]),
                .reg45        (o_d_reg[16][45]),
                .reg46        (o_d_reg[16][46]),
                .reg47        (o_d_reg[16][47]),
                .reg48        (o_d_reg[16][48]),
                .reg49        (o_d_reg[16][49]),
                .reg50        (o_d_reg[16][50]),
                .reg51        (o_d_reg[16][51]),
                .reg52        (o_d_reg[16][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf17
        (
                .din        (o_d_rowBuf[16]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[17]),
                .reg01        (o_d_reg[17][1]),
                .reg02        (o_d_reg[17][2]),
                .reg03        (o_d_reg[17][3]),
                .reg04        (o_d_reg[17][4]),
                .reg05        (o_d_reg[17][5]),
                .reg06        (o_d_reg[17][6]),
                .reg07        (o_d_reg[17][7]),
                .reg08        (o_d_reg[17][8]),
                .reg09        (o_d_reg[17][9]),
                .reg10        (o_d_reg[17][10]),
                .reg11        (o_d_reg[17][11]),
                .reg12        (o_d_reg[17][12]),
                .reg13        (o_d_reg[17][13]),
                .reg14        (o_d_reg[17][14]),
                .reg15        (o_d_reg[17][15]),
                .reg16        (o_d_reg[17][16]),
                .reg17        (o_d_reg[17][17]),
                .reg18        (o_d_reg[17][18]),
                .reg19        (o_d_reg[17][19]),
                .reg20        (o_d_reg[17][20]),
                .reg21        (o_d_reg[17][21]),
                .reg22        (o_d_reg[17][22]),
                .reg23        (o_d_reg[17][23]),
                .reg24        (o_d_reg[17][24]),
                .reg25        (o_d_reg[17][25]),
                .reg26        (o_d_reg[17][26]),
                .reg27        (o_d_reg[17][27]),
                .reg28        (o_d_reg[17][28]),
                .reg29        (o_d_reg[17][29]),
                .reg30        (o_d_reg[17][30]),
                .reg31        (o_d_reg[17][31]),
                .reg32        (o_d_reg[17][32]),
                .reg33        (o_d_reg[17][33]),
                .reg34        (o_d_reg[17][34]),
                .reg35        (o_d_reg[17][35]),
                .reg36        (o_d_reg[17][36]),
                .reg37        (o_d_reg[17][37]),
                .reg38        (o_d_reg[17][38]),
                .reg39        (o_d_reg[17][39]),
                .reg40        (o_d_reg[17][40]),
                .reg41        (o_d_reg[17][41]),
                .reg42        (o_d_reg[17][42]),
                .reg43        (o_d_reg[17][43]),
                .reg44        (o_d_reg[17][44]),
                .reg45        (o_d_reg[17][45]),
                .reg46        (o_d_reg[17][46]),
                .reg47        (o_d_reg[17][47]),
                .reg48        (o_d_reg[17][48]),
                .reg49        (o_d_reg[17][49]),
                .reg50        (o_d_reg[17][50]),
                .reg51        (o_d_reg[17][51]),
                .reg52        (o_d_reg[17][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf18
        (
                .din        (o_d_rowBuf[17]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[18]),
                .reg01        (o_d_reg[18][1]),
                .reg02        (o_d_reg[18][2]),
                .reg03        (o_d_reg[18][3]),
                .reg04        (o_d_reg[18][4]),
                .reg05        (o_d_reg[18][5]),
                .reg06        (o_d_reg[18][6]),
                .reg07        (o_d_reg[18][7]),
                .reg08        (o_d_reg[18][8]),
                .reg09        (o_d_reg[18][9]),
                .reg10        (o_d_reg[18][10]),
                .reg11        (o_d_reg[18][11]),
                .reg12        (o_d_reg[18][12]),
                .reg13        (o_d_reg[18][13]),
                .reg14        (o_d_reg[18][14]),
                .reg15        (o_d_reg[18][15]),
                .reg16        (o_d_reg[18][16]),
                .reg17        (o_d_reg[18][17]),
                .reg18        (o_d_reg[18][18]),
                .reg19        (o_d_reg[18][19]),
                .reg20        (o_d_reg[18][20]),
                .reg21        (o_d_reg[18][21]),
                .reg22        (o_d_reg[18][22]),
                .reg23        (o_d_reg[18][23]),
                .reg24        (o_d_reg[18][24]),
                .reg25        (o_d_reg[18][25]),
                .reg26        (o_d_reg[18][26]),
                .reg27        (o_d_reg[18][27]),
                .reg28        (o_d_reg[18][28]),
                .reg29        (o_d_reg[18][29]),
                .reg30        (o_d_reg[18][30]),
                .reg31        (o_d_reg[18][31]),
                .reg32        (o_d_reg[18][32]),
                .reg33        (o_d_reg[18][33]),
                .reg34        (o_d_reg[18][34]),
                .reg35        (o_d_reg[18][35]),
                .reg36        (o_d_reg[18][36]),
                .reg37        (o_d_reg[18][37]),
                .reg38        (o_d_reg[18][38]),
                .reg39        (o_d_reg[18][39]),
                .reg40        (o_d_reg[18][40]),
                .reg41        (o_d_reg[18][41]),
                .reg42        (o_d_reg[18][42]),
                .reg43        (o_d_reg[18][43]),
                .reg44        (o_d_reg[18][44]),
                .reg45        (o_d_reg[18][45]),
                .reg46        (o_d_reg[18][46]),
                .reg47        (o_d_reg[18][47]),
                .reg48        (o_d_reg[18][48]),
                .reg49        (o_d_reg[18][49]),
                .reg50        (o_d_reg[18][50]),
                .reg51        (o_d_reg[18][51]),
                .reg52        (o_d_reg[18][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf19
        (
                .din        (o_d_rowBuf[18]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[19]),
                .reg01        (o_d_reg[19][1]),
                .reg02        (o_d_reg[19][2]),
                .reg03        (o_d_reg[19][3]),
                .reg04        (o_d_reg[19][4]),
                .reg05        (o_d_reg[19][5]),
                .reg06        (o_d_reg[19][6]),
                .reg07        (o_d_reg[19][7]),
                .reg08        (o_d_reg[19][8]),
                .reg09        (o_d_reg[19][9]),
                .reg10        (o_d_reg[19][10]),
                .reg11        (o_d_reg[19][11]),
                .reg12        (o_d_reg[19][12]),
                .reg13        (o_d_reg[19][13]),
                .reg14        (o_d_reg[19][14]),
                .reg15        (o_d_reg[19][15]),
                .reg16        (o_d_reg[19][16]),
                .reg17        (o_d_reg[19][17]),
                .reg18        (o_d_reg[19][18]),
                .reg19        (o_d_reg[19][19]),
                .reg20        (o_d_reg[19][20]),
                .reg21        (o_d_reg[19][21]),
                .reg22        (o_d_reg[19][22]),
                .reg23        (o_d_reg[19][23]),
                .reg24        (o_d_reg[19][24]),
                .reg25        (o_d_reg[19][25]),
                .reg26        (o_d_reg[19][26]),
                .reg27        (o_d_reg[19][27]),
                .reg28        (o_d_reg[19][28]),
                .reg29        (o_d_reg[19][29]),
                .reg30        (o_d_reg[19][30]),
                .reg31        (o_d_reg[19][31]),
                .reg32        (o_d_reg[19][32]),
                .reg33        (o_d_reg[19][33]),
                .reg34        (o_d_reg[19][34]),
                .reg35        (o_d_reg[19][35]),
                .reg36        (o_d_reg[19][36]),
                .reg37        (o_d_reg[19][37]),
                .reg38        (o_d_reg[19][38]),
                .reg39        (o_d_reg[19][39]),
                .reg40        (o_d_reg[19][40]),
                .reg41        (o_d_reg[19][41]),
                .reg42        (o_d_reg[19][42]),
                .reg43        (o_d_reg[19][43]),
                .reg44        (o_d_reg[19][44]),
                .reg45        (o_d_reg[19][45]),
                .reg46        (o_d_reg[19][46]),
                .reg47        (o_d_reg[19][47]),
                .reg48        (o_d_reg[19][48]),
                .reg49        (o_d_reg[19][49]),
                .reg50        (o_d_reg[19][50]),
                .reg51        (o_d_reg[19][51]),
                .reg52        (o_d_reg[19][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf20
        (
                .din        (o_d_rowBuf[19]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[20]),
                .reg01        (o_d_reg[20][1]),
                .reg02        (o_d_reg[20][2]),
                .reg03        (o_d_reg[20][3]),
                .reg04        (o_d_reg[20][4]),
                .reg05        (o_d_reg[20][5]),
                .reg06        (o_d_reg[20][6]),
                .reg07        (o_d_reg[20][7]),
                .reg08        (o_d_reg[20][8]),
                .reg09        (o_d_reg[20][9]),
                .reg10        (o_d_reg[20][10]),
                .reg11        (o_d_reg[20][11]),
                .reg12        (o_d_reg[20][12]),
                .reg13        (o_d_reg[20][13]),
                .reg14        (o_d_reg[20][14]),
                .reg15        (o_d_reg[20][15]),
                .reg16        (o_d_reg[20][16]),
                .reg17        (o_d_reg[20][17]),
                .reg18        (o_d_reg[20][18]),
                .reg19        (o_d_reg[20][19]),
                .reg20        (o_d_reg[20][20]),
                .reg21        (o_d_reg[20][21]),
                .reg22        (o_d_reg[20][22]),
                .reg23        (o_d_reg[20][23]),
                .reg24        (o_d_reg[20][24]),
                .reg25        (o_d_reg[20][25]),
                .reg26        (o_d_reg[20][26]),
                .reg27        (o_d_reg[20][27]),
                .reg28        (o_d_reg[20][28]),
                .reg29        (o_d_reg[20][29]),
                .reg30        (o_d_reg[20][30]),
                .reg31        (o_d_reg[20][31]),
                .reg32        (o_d_reg[20][32]),
                .reg33        (o_d_reg[20][33]),
                .reg34        (o_d_reg[20][34]),
                .reg35        (o_d_reg[20][35]),
                .reg36        (o_d_reg[20][36]),
                .reg37        (o_d_reg[20][37]),
                .reg38        (o_d_reg[20][38]),
                .reg39        (o_d_reg[20][39]),
                .reg40        (o_d_reg[20][40]),
                .reg41        (o_d_reg[20][41]),
                .reg42        (o_d_reg[20][42]),
                .reg43        (o_d_reg[20][43]),
                .reg44        (o_d_reg[20][44]),
                .reg45        (o_d_reg[20][45]),
                .reg46        (o_d_reg[20][46]),
                .reg47        (o_d_reg[20][47]),
                .reg48        (o_d_reg[20][48]),
                .reg49        (o_d_reg[20][49]),
                .reg50        (o_d_reg[20][50]),
                .reg51        (o_d_reg[20][51]),
                .reg52        (o_d_reg[20][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf21
        (
                .din        (o_d_rowBuf[20]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[21]),
                .reg01        (o_d_reg[21][1]),
                .reg02        (o_d_reg[21][2]),
                .reg03        (o_d_reg[21][3]),
                .reg04        (o_d_reg[21][4]),
                .reg05        (o_d_reg[21][5]),
                .reg06        (o_d_reg[21][6]),
                .reg07        (o_d_reg[21][7]),
                .reg08        (o_d_reg[21][8]),
                .reg09        (o_d_reg[21][9]),
                .reg10        (o_d_reg[21][10]),
                .reg11        (o_d_reg[21][11]),
                .reg12        (o_d_reg[21][12]),
                .reg13        (o_d_reg[21][13]),
                .reg14        (o_d_reg[21][14]),
                .reg15        (o_d_reg[21][15]),
                .reg16        (o_d_reg[21][16]),
                .reg17        (o_d_reg[21][17]),
                .reg18        (o_d_reg[21][18]),
                .reg19        (o_d_reg[21][19]),
                .reg20        (o_d_reg[21][20]),
                .reg21        (o_d_reg[21][21]),
                .reg22        (o_d_reg[21][22]),
                .reg23        (o_d_reg[21][23]),
                .reg24        (o_d_reg[21][24]),
                .reg25        (o_d_reg[21][25]),
                .reg26        (o_d_reg[21][26]),
                .reg27        (o_d_reg[21][27]),
                .reg28        (o_d_reg[21][28]),
                .reg29        (o_d_reg[21][29]),
                .reg30        (o_d_reg[21][30]),
                .reg31        (o_d_reg[21][31]),
                .reg32        (o_d_reg[21][32]),
                .reg33        (o_d_reg[21][33]),
                .reg34        (o_d_reg[21][34]),
                .reg35        (o_d_reg[21][35]),
                .reg36        (o_d_reg[21][36]),
                .reg37        (o_d_reg[21][37]),
                .reg38        (o_d_reg[21][38]),
                .reg39        (o_d_reg[21][39]),
                .reg40        (o_d_reg[21][40]),
                .reg41        (o_d_reg[21][41]),
                .reg42        (o_d_reg[21][42]),
                .reg43        (o_d_reg[21][43]),
                .reg44        (o_d_reg[21][44]),
                .reg45        (o_d_reg[21][45]),
                .reg46        (o_d_reg[21][46]),
                .reg47        (o_d_reg[21][47]),
                .reg48        (o_d_reg[21][48]),
                .reg49        (o_d_reg[21][49]),
                .reg50        (o_d_reg[21][50]),
                .reg51        (o_d_reg[21][51]),
                .reg52        (o_d_reg[21][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf22
        (
                .din        (o_d_rowBuf[21]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[22]),
                .reg01        (o_d_reg[22][1]),
                .reg02        (o_d_reg[22][2]),
                .reg03        (o_d_reg[22][3]),
                .reg04        (o_d_reg[22][4]),
                .reg05        (o_d_reg[22][5]),
                .reg06        (o_d_reg[22][6]),
                .reg07        (o_d_reg[22][7]),
                .reg08        (o_d_reg[22][8]),
                .reg09        (o_d_reg[22][9]),
                .reg10        (o_d_reg[22][10]),
                .reg11        (o_d_reg[22][11]),
                .reg12        (o_d_reg[22][12]),
                .reg13        (o_d_reg[22][13]),
                .reg14        (o_d_reg[22][14]),
                .reg15        (o_d_reg[22][15]),
                .reg16        (o_d_reg[22][16]),
                .reg17        (o_d_reg[22][17]),
                .reg18        (o_d_reg[22][18]),
                .reg19        (o_d_reg[22][19]),
                .reg20        (o_d_reg[22][20]),
                .reg21        (o_d_reg[22][21]),
                .reg22        (o_d_reg[22][22]),
                .reg23        (o_d_reg[22][23]),
                .reg24        (o_d_reg[22][24]),
                .reg25        (o_d_reg[22][25]),
                .reg26        (o_d_reg[22][26]),
                .reg27        (o_d_reg[22][27]),
                .reg28        (o_d_reg[22][28]),
                .reg29        (o_d_reg[22][29]),
                .reg30        (o_d_reg[22][30]),
                .reg31        (o_d_reg[22][31]),
                .reg32        (o_d_reg[22][32]),
                .reg33        (o_d_reg[22][33]),
                .reg34        (o_d_reg[22][34]),
                .reg35        (o_d_reg[22][35]),
                .reg36        (o_d_reg[22][36]),
                .reg37        (o_d_reg[22][37]),
                .reg38        (o_d_reg[22][38]),
                .reg39        (o_d_reg[22][39]),
                .reg40        (o_d_reg[22][40]),
                .reg41        (o_d_reg[22][41]),
                .reg42        (o_d_reg[22][42]),
                .reg43        (o_d_reg[22][43]),
                .reg44        (o_d_reg[22][44]),
                .reg45        (o_d_reg[22][45]),
                .reg46        (o_d_reg[22][46]),
                .reg47        (o_d_reg[22][47]),
                .reg48        (o_d_reg[22][48]),
                .reg49        (o_d_reg[22][49]),
                .reg50        (o_d_reg[22][50]),
                .reg51        (o_d_reg[22][51]),
                .reg52        (o_d_reg[22][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf23
        (
                .din        (o_d_rowBuf[22]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[23]),
                .reg01        (o_d_reg[23][1]),
                .reg02        (o_d_reg[23][2]),
                .reg03        (o_d_reg[23][3]),
                .reg04        (o_d_reg[23][4]),
                .reg05        (o_d_reg[23][5]),
                .reg06        (o_d_reg[23][6]),
                .reg07        (o_d_reg[23][7]),
                .reg08        (o_d_reg[23][8]),
                .reg09        (o_d_reg[23][9]),
                .reg10        (o_d_reg[23][10]),
                .reg11        (o_d_reg[23][11]),
                .reg12        (o_d_reg[23][12]),
                .reg13        (o_d_reg[23][13]),
                .reg14        (o_d_reg[23][14]),
                .reg15        (o_d_reg[23][15]),
                .reg16        (o_d_reg[23][16]),
                .reg17        (o_d_reg[23][17]),
                .reg18        (o_d_reg[23][18]),
                .reg19        (o_d_reg[23][19]),
                .reg20        (o_d_reg[23][20]),
                .reg21        (o_d_reg[23][21]),
                .reg22        (o_d_reg[23][22]),
                .reg23        (o_d_reg[23][23]),
                .reg24        (o_d_reg[23][24]),
                .reg25        (o_d_reg[23][25]),
                .reg26        (o_d_reg[23][26]),
                .reg27        (o_d_reg[23][27]),
                .reg28        (o_d_reg[23][28]),
                .reg29        (o_d_reg[23][29]),
                .reg30        (o_d_reg[23][30]),
                .reg31        (o_d_reg[23][31]),
                .reg32        (o_d_reg[23][32]),
                .reg33        (o_d_reg[23][33]),
                .reg34        (o_d_reg[23][34]),
                .reg35        (o_d_reg[23][35]),
                .reg36        (o_d_reg[23][36]),
                .reg37        (o_d_reg[23][37]),
                .reg38        (o_d_reg[23][38]),
                .reg39        (o_d_reg[23][39]),
                .reg40        (o_d_reg[23][40]),
                .reg41        (o_d_reg[23][41]),
                .reg42        (o_d_reg[23][42]),
                .reg43        (o_d_reg[23][43]),
                .reg44        (o_d_reg[23][44]),
                .reg45        (o_d_reg[23][45]),
                .reg46        (o_d_reg[23][46]),
                .reg47        (o_d_reg[23][47]),
                .reg48        (o_d_reg[23][48]),
                .reg49        (o_d_reg[23][49]),
                .reg50        (o_d_reg[23][50]),
                .reg51        (o_d_reg[23][51]),
                .reg52        (o_d_reg[23][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf24
        (
                .din        (o_d_rowBuf[23]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[24]),
                .reg01        (o_d_reg[24][1]),
                .reg02        (o_d_reg[24][2]),
                .reg03        (o_d_reg[24][3]),
                .reg04        (o_d_reg[24][4]),
                .reg05        (o_d_reg[24][5]),
                .reg06        (o_d_reg[24][6]),
                .reg07        (o_d_reg[24][7]),
                .reg08        (o_d_reg[24][8]),
                .reg09        (o_d_reg[24][9]),
                .reg10        (o_d_reg[24][10]),
                .reg11        (o_d_reg[24][11]),
                .reg12        (o_d_reg[24][12]),
                .reg13        (o_d_reg[24][13]),
                .reg14        (o_d_reg[24][14]),
                .reg15        (o_d_reg[24][15]),
                .reg16        (o_d_reg[24][16]),
                .reg17        (o_d_reg[24][17]),
                .reg18        (o_d_reg[24][18]),
                .reg19        (o_d_reg[24][19]),
                .reg20        (o_d_reg[24][20]),
                .reg21        (o_d_reg[24][21]),
                .reg22        (o_d_reg[24][22]),
                .reg23        (o_d_reg[24][23]),
                .reg24        (o_d_reg[24][24]),
                .reg25        (o_d_reg[24][25]),
                .reg26        (o_d_reg[24][26]),
                .reg27        (o_d_reg[24][27]),
                .reg28        (o_d_reg[24][28]),
                .reg29        (o_d_reg[24][29]),
                .reg30        (o_d_reg[24][30]),
                .reg31        (o_d_reg[24][31]),
                .reg32        (o_d_reg[24][32]),
                .reg33        (o_d_reg[24][33]),
                .reg34        (o_d_reg[24][34]),
                .reg35        (o_d_reg[24][35]),
                .reg36        (o_d_reg[24][36]),
                .reg37        (o_d_reg[24][37]),
                .reg38        (o_d_reg[24][38]),
                .reg39        (o_d_reg[24][39]),
                .reg40        (o_d_reg[24][40]),
                .reg41        (o_d_reg[24][41]),
                .reg42        (o_d_reg[24][42]),
                .reg43        (o_d_reg[24][43]),
                .reg44        (o_d_reg[24][44]),
                .reg45        (o_d_reg[24][45]),
                .reg46        (o_d_reg[24][46]),
                .reg47        (o_d_reg[24][47]),
                .reg48        (o_d_reg[24][48]),
                .reg49        (o_d_reg[24][49]),
                .reg50        (o_d_reg[24][50]),
                .reg51        (o_d_reg[24][51]),
                .reg52        (o_d_reg[24][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf25
        (
                .din        (o_d_rowBuf[24]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[25]),
                .reg01        (o_d_reg[25][1]),
                .reg02        (o_d_reg[25][2]),
                .reg03        (o_d_reg[25][3]),
                .reg04        (o_d_reg[25][4]),
                .reg05        (o_d_reg[25][5]),
                .reg06        (o_d_reg[25][6]),
                .reg07        (o_d_reg[25][7]),
                .reg08        (o_d_reg[25][8]),
                .reg09        (o_d_reg[25][9]),
                .reg10        (o_d_reg[25][10]),
                .reg11        (o_d_reg[25][11]),
                .reg12        (o_d_reg[25][12]),
                .reg13        (o_d_reg[25][13]),
                .reg14        (o_d_reg[25][14]),
                .reg15        (o_d_reg[25][15]),
                .reg16        (o_d_reg[25][16]),
                .reg17        (o_d_reg[25][17]),
                .reg18        (o_d_reg[25][18]),
                .reg19        (o_d_reg[25][19]),
                .reg20        (o_d_reg[25][20]),
                .reg21        (o_d_reg[25][21]),
                .reg22        (o_d_reg[25][22]),
                .reg23        (o_d_reg[25][23]),
                .reg24        (o_d_reg[25][24]),
                .reg25        (o_d_reg[25][25]),
                .reg26        (o_d_reg[25][26]),
                .reg27        (o_d_reg[25][27]),
                .reg28        (o_d_reg[25][28]),
                .reg29        (o_d_reg[25][29]),
                .reg30        (o_d_reg[25][30]),
                .reg31        (o_d_reg[25][31]),
                .reg32        (o_d_reg[25][32]),
                .reg33        (o_d_reg[25][33]),
                .reg34        (o_d_reg[25][34]),
                .reg35        (o_d_reg[25][35]),
                .reg36        (o_d_reg[25][36]),
                .reg37        (o_d_reg[25][37]),
                .reg38        (o_d_reg[25][38]),
                .reg39        (o_d_reg[25][39]),
                .reg40        (o_d_reg[25][40]),
                .reg41        (o_d_reg[25][41]),
                .reg42        (o_d_reg[25][42]),
                .reg43        (o_d_reg[25][43]),
                .reg44        (o_d_reg[25][44]),
                .reg45        (o_d_reg[25][45]),
                .reg46        (o_d_reg[25][46]),
                .reg47        (o_d_reg[25][47]),
                .reg48        (o_d_reg[25][48]),
                .reg49        (o_d_reg[25][49]),
                .reg50        (o_d_reg[25][50]),
                .reg51        (o_d_reg[25][51]),
                .reg52        (o_d_reg[25][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf26
        (
                .din        (o_d_rowBuf[25]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[26]),
                .reg01        (o_d_reg[26][1]),
                .reg02        (o_d_reg[26][2]),
                .reg03        (o_d_reg[26][3]),
                .reg04        (o_d_reg[26][4]),
                .reg05        (o_d_reg[26][5]),
                .reg06        (o_d_reg[26][6]),
                .reg07        (o_d_reg[26][7]),
                .reg08        (o_d_reg[26][8]),
                .reg09        (o_d_reg[26][9]),
                .reg10        (o_d_reg[26][10]),
                .reg11        (o_d_reg[26][11]),
                .reg12        (o_d_reg[26][12]),
                .reg13        (o_d_reg[26][13]),
                .reg14        (o_d_reg[26][14]),
                .reg15        (o_d_reg[26][15]),
                .reg16        (o_d_reg[26][16]),
                .reg17        (o_d_reg[26][17]),
                .reg18        (o_d_reg[26][18]),
                .reg19        (o_d_reg[26][19]),
                .reg20        (o_d_reg[26][20]),
                .reg21        (o_d_reg[26][21]),
                .reg22        (o_d_reg[26][22]),
                .reg23        (o_d_reg[26][23]),
                .reg24        (o_d_reg[26][24]),
                .reg25        (o_d_reg[26][25]),
                .reg26        (o_d_reg[26][26]),
                .reg27        (o_d_reg[26][27]),
                .reg28        (o_d_reg[26][28]),
                .reg29        (o_d_reg[26][29]),
                .reg30        (o_d_reg[26][30]),
                .reg31        (o_d_reg[26][31]),
                .reg32        (o_d_reg[26][32]),
                .reg33        (o_d_reg[26][33]),
                .reg34        (o_d_reg[26][34]),
                .reg35        (o_d_reg[26][35]),
                .reg36        (o_d_reg[26][36]),
                .reg37        (o_d_reg[26][37]),
                .reg38        (o_d_reg[26][38]),
                .reg39        (o_d_reg[26][39]),
                .reg40        (o_d_reg[26][40]),
                .reg41        (o_d_reg[26][41]),
                .reg42        (o_d_reg[26][42]),
                .reg43        (o_d_reg[26][43]),
                .reg44        (o_d_reg[26][44]),
                .reg45        (o_d_reg[26][45]),
                .reg46        (o_d_reg[26][46]),
                .reg47        (o_d_reg[26][47]),
                .reg48        (o_d_reg[26][48]),
                .reg49        (o_d_reg[26][49]),
                .reg50        (o_d_reg[26][50]),
                .reg51        (o_d_reg[26][51]),
                .reg52        (o_d_reg[26][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf27
        (
                .din        (o_d_rowBuf[26]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[27]),
                .reg01        (o_d_reg[27][1]),
                .reg02        (o_d_reg[27][2]),
                .reg03        (o_d_reg[27][3]),
                .reg04        (o_d_reg[27][4]),
                .reg05        (o_d_reg[27][5]),
                .reg06        (o_d_reg[27][6]),
                .reg07        (o_d_reg[27][7]),
                .reg08        (o_d_reg[27][8]),
                .reg09        (o_d_reg[27][9]),
                .reg10        (o_d_reg[27][10]),
                .reg11        (o_d_reg[27][11]),
                .reg12        (o_d_reg[27][12]),
                .reg13        (o_d_reg[27][13]),
                .reg14        (o_d_reg[27][14]),
                .reg15        (o_d_reg[27][15]),
                .reg16        (o_d_reg[27][16]),
                .reg17        (o_d_reg[27][17]),
                .reg18        (o_d_reg[27][18]),
                .reg19        (o_d_reg[27][19]),
                .reg20        (o_d_reg[27][20]),
                .reg21        (o_d_reg[27][21]),
                .reg22        (o_d_reg[27][22]),
                .reg23        (o_d_reg[27][23]),
                .reg24        (o_d_reg[27][24]),
                .reg25        (o_d_reg[27][25]),
                .reg26        (o_d_reg[27][26]),
                .reg27        (o_d_reg[27][27]),
                .reg28        (o_d_reg[27][28]),
                .reg29        (o_d_reg[27][29]),
                .reg30        (o_d_reg[27][30]),
                .reg31        (o_d_reg[27][31]),
                .reg32        (o_d_reg[27][32]),
                .reg33        (o_d_reg[27][33]),
                .reg34        (o_d_reg[27][34]),
                .reg35        (o_d_reg[27][35]),
                .reg36        (o_d_reg[27][36]),
                .reg37        (o_d_reg[27][37]),
                .reg38        (o_d_reg[27][38]),
                .reg39        (o_d_reg[27][39]),
                .reg40        (o_d_reg[27][40]),
                .reg41        (o_d_reg[27][41]),
                .reg42        (o_d_reg[27][42]),
                .reg43        (o_d_reg[27][43]),
                .reg44        (o_d_reg[27][44]),
                .reg45        (o_d_reg[27][45]),
                .reg46        (o_d_reg[27][46]),
                .reg47        (o_d_reg[27][47]),
                .reg48        (o_d_reg[27][48]),
                .reg49        (o_d_reg[27][49]),
                .reg50        (o_d_reg[27][50]),
                .reg51        (o_d_reg[27][51]),
                .reg52        (o_d_reg[27][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf28
        (
                .din        (o_d_rowBuf[27]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[28]),
                .reg01        (o_d_reg[28][1]),
                .reg02        (o_d_reg[28][2]),
                .reg03        (o_d_reg[28][3]),
                .reg04        (o_d_reg[28][4]),
                .reg05        (o_d_reg[28][5]),
                .reg06        (o_d_reg[28][6]),
                .reg07        (o_d_reg[28][7]),
                .reg08        (o_d_reg[28][8]),
                .reg09        (o_d_reg[28][9]),
                .reg10        (o_d_reg[28][10]),
                .reg11        (o_d_reg[28][11]),
                .reg12        (o_d_reg[28][12]),
                .reg13        (o_d_reg[28][13]),
                .reg14        (o_d_reg[28][14]),
                .reg15        (o_d_reg[28][15]),
                .reg16        (o_d_reg[28][16]),
                .reg17        (o_d_reg[28][17]),
                .reg18        (o_d_reg[28][18]),
                .reg19        (o_d_reg[28][19]),
                .reg20        (o_d_reg[28][20]),
                .reg21        (o_d_reg[28][21]),
                .reg22        (o_d_reg[28][22]),
                .reg23        (o_d_reg[28][23]),
                .reg24        (o_d_reg[28][24]),
                .reg25        (o_d_reg[28][25]),
                .reg26        (o_d_reg[28][26]),
                .reg27        (o_d_reg[28][27]),
                .reg28        (o_d_reg[28][28]),
                .reg29        (o_d_reg[28][29]),
                .reg30        (o_d_reg[28][30]),
                .reg31        (o_d_reg[28][31]),
                .reg32        (o_d_reg[28][32]),
                .reg33        (o_d_reg[28][33]),
                .reg34        (o_d_reg[28][34]),
                .reg35        (o_d_reg[28][35]),
                .reg36        (o_d_reg[28][36]),
                .reg37        (o_d_reg[28][37]),
                .reg38        (o_d_reg[28][38]),
                .reg39        (o_d_reg[28][39]),
                .reg40        (o_d_reg[28][40]),
                .reg41        (o_d_reg[28][41]),
                .reg42        (o_d_reg[28][42]),
                .reg43        (o_d_reg[28][43]),
                .reg44        (o_d_reg[28][44]),
                .reg45        (o_d_reg[28][45]),
                .reg46        (o_d_reg[28][46]),
                .reg47        (o_d_reg[28][47]),
                .reg48        (o_d_reg[28][48]),
                .reg49        (o_d_reg[28][49]),
                .reg50        (o_d_reg[28][50]),
                .reg51        (o_d_reg[28][51]),
                .reg52        (o_d_reg[28][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf29
        (
                .din        (o_d_rowBuf[28]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[29]),
                .reg01        (o_d_reg[29][1]),
                .reg02        (o_d_reg[29][2]),
                .reg03        (o_d_reg[29][3]),
                .reg04        (o_d_reg[29][4]),
                .reg05        (o_d_reg[29][5]),
                .reg06        (o_d_reg[29][6]),
                .reg07        (o_d_reg[29][7]),
                .reg08        (o_d_reg[29][8]),
                .reg09        (o_d_reg[29][9]),
                .reg10        (o_d_reg[29][10]),
                .reg11        (o_d_reg[29][11]),
                .reg12        (o_d_reg[29][12]),
                .reg13        (o_d_reg[29][13]),
                .reg14        (o_d_reg[29][14]),
                .reg15        (o_d_reg[29][15]),
                .reg16        (o_d_reg[29][16]),
                .reg17        (o_d_reg[29][17]),
                .reg18        (o_d_reg[29][18]),
                .reg19        (o_d_reg[29][19]),
                .reg20        (o_d_reg[29][20]),
                .reg21        (o_d_reg[29][21]),
                .reg22        (o_d_reg[29][22]),
                .reg23        (o_d_reg[29][23]),
                .reg24        (o_d_reg[29][24]),
                .reg25        (o_d_reg[29][25]),
                .reg26        (o_d_reg[29][26]),
                .reg27        (o_d_reg[29][27]),
                .reg28        (o_d_reg[29][28]),
                .reg29        (o_d_reg[29][29]),
                .reg30        (o_d_reg[29][30]),
                .reg31        (o_d_reg[29][31]),
                .reg32        (o_d_reg[29][32]),
                .reg33        (o_d_reg[29][33]),
                .reg34        (o_d_reg[29][34]),
                .reg35        (o_d_reg[29][35]),
                .reg36        (o_d_reg[29][36]),
                .reg37        (o_d_reg[29][37]),
                .reg38        (o_d_reg[29][38]),
                .reg39        (o_d_reg[29][39]),
                .reg40        (o_d_reg[29][40]),
                .reg41        (o_d_reg[29][41]),
                .reg42        (o_d_reg[29][42]),
                .reg43        (o_d_reg[29][43]),
                .reg44        (o_d_reg[29][44]),
                .reg45        (o_d_reg[29][45]),
                .reg46        (o_d_reg[29][46]),
                .reg47        (o_d_reg[29][47]),
                .reg48        (o_d_reg[29][48]),
                .reg49        (o_d_reg[29][49]),
                .reg50        (o_d_reg[29][50]),
                .reg51        (o_d_reg[29][51]),
                .reg52        (o_d_reg[29][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf30
        (
                .din        (o_d_rowBuf[29]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[30]),
                .reg01        (o_d_reg[30][1]),
                .reg02        (o_d_reg[30][2]),
                .reg03        (o_d_reg[30][3]),
                .reg04        (o_d_reg[30][4]),
                .reg05        (o_d_reg[30][5]),
                .reg06        (o_d_reg[30][6]),
                .reg07        (o_d_reg[30][7]),
                .reg08        (o_d_reg[30][8]),
                .reg09        (o_d_reg[30][9]),
                .reg10        (o_d_reg[30][10]),
                .reg11        (o_d_reg[30][11]),
                .reg12        (o_d_reg[30][12]),
                .reg13        (o_d_reg[30][13]),
                .reg14        (o_d_reg[30][14]),
                .reg15        (o_d_reg[30][15]),
                .reg16        (o_d_reg[30][16]),
                .reg17        (o_d_reg[30][17]),
                .reg18        (o_d_reg[30][18]),
                .reg19        (o_d_reg[30][19]),
                .reg20        (o_d_reg[30][20]),
                .reg21        (o_d_reg[30][21]),
                .reg22        (o_d_reg[30][22]),
                .reg23        (o_d_reg[30][23]),
                .reg24        (o_d_reg[30][24]),
                .reg25        (o_d_reg[30][25]),
                .reg26        (o_d_reg[30][26]),
                .reg27        (o_d_reg[30][27]),
                .reg28        (o_d_reg[30][28]),
                .reg29        (o_d_reg[30][29]),
                .reg30        (o_d_reg[30][30]),
                .reg31        (o_d_reg[30][31]),
                .reg32        (o_d_reg[30][32]),
                .reg33        (o_d_reg[30][33]),
                .reg34        (o_d_reg[30][34]),
                .reg35        (o_d_reg[30][35]),
                .reg36        (o_d_reg[30][36]),
                .reg37        (o_d_reg[30][37]),
                .reg38        (o_d_reg[30][38]),
                .reg39        (o_d_reg[30][39]),
                .reg40        (o_d_reg[30][40]),
                .reg41        (o_d_reg[30][41]),
                .reg42        (o_d_reg[30][42]),
                .reg43        (o_d_reg[30][43]),
                .reg44        (o_d_reg[30][44]),
                .reg45        (o_d_reg[30][45]),
                .reg46        (o_d_reg[30][46]),
                .reg47        (o_d_reg[30][47]),
                .reg48        (o_d_reg[30][48]),
                .reg49        (o_d_reg[30][49]),
                .reg50        (o_d_reg[30][50]),
                .reg51        (o_d_reg[30][51]),
                .reg52        (o_d_reg[30][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf31
        (
                .din        (o_d_rowBuf[30]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[31]),
                .reg01        (o_d_reg[31][1]),
                .reg02        (o_d_reg[31][2]),
                .reg03        (o_d_reg[31][3]),
                .reg04        (o_d_reg[31][4]),
                .reg05        (o_d_reg[31][5]),
                .reg06        (o_d_reg[31][6]),
                .reg07        (o_d_reg[31][7]),
                .reg08        (o_d_reg[31][8]),
                .reg09        (o_d_reg[31][9]),
                .reg10        (o_d_reg[31][10]),
                .reg11        (o_d_reg[31][11]),
                .reg12        (o_d_reg[31][12]),
                .reg13        (o_d_reg[31][13]),
                .reg14        (o_d_reg[31][14]),
                .reg15        (o_d_reg[31][15]),
                .reg16        (o_d_reg[31][16]),
                .reg17        (o_d_reg[31][17]),
                .reg18        (o_d_reg[31][18]),
                .reg19        (o_d_reg[31][19]),
                .reg20        (o_d_reg[31][20]),
                .reg21        (o_d_reg[31][21]),
                .reg22        (o_d_reg[31][22]),
                .reg23        (o_d_reg[31][23]),
                .reg24        (o_d_reg[31][24]),
                .reg25        (o_d_reg[31][25]),
                .reg26        (o_d_reg[31][26]),
                .reg27        (o_d_reg[31][27]),
                .reg28        (o_d_reg[31][28]),
                .reg29        (o_d_reg[31][29]),
                .reg30        (o_d_reg[31][30]),
                .reg31        (o_d_reg[31][31]),
                .reg32        (o_d_reg[31][32]),
                .reg33        (o_d_reg[31][33]),
                .reg34        (o_d_reg[31][34]),
                .reg35        (o_d_reg[31][35]),
                .reg36        (o_d_reg[31][36]),
                .reg37        (o_d_reg[31][37]),
                .reg38        (o_d_reg[31][38]),
                .reg39        (o_d_reg[31][39]),
                .reg40        (o_d_reg[31][40]),
                .reg41        (o_d_reg[31][41]),
                .reg42        (o_d_reg[31][42]),
                .reg43        (o_d_reg[31][43]),
                .reg44        (o_d_reg[31][44]),
                .reg45        (o_d_reg[31][45]),
                .reg46        (o_d_reg[31][46]),
                .reg47        (o_d_reg[31][47]),
                .reg48        (o_d_reg[31][48]),
                .reg49        (o_d_reg[31][49]),
                .reg50        (o_d_reg[31][50]),
                .reg51        (o_d_reg[31][51]),
                .reg52        (o_d_reg[31][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf32
        (
                .din        (o_d_rowBuf[31]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[32]),
                .reg01        (o_d_reg[32][1]),
                .reg02        (o_d_reg[32][2]),
                .reg03        (o_d_reg[32][3]),
                .reg04        (o_d_reg[32][4]),
                .reg05        (o_d_reg[32][5]),
                .reg06        (o_d_reg[32][6]),
                .reg07        (o_d_reg[32][7]),
                .reg08        (o_d_reg[32][8]),
                .reg09        (o_d_reg[32][9]),
                .reg10        (o_d_reg[32][10]),
                .reg11        (o_d_reg[32][11]),
                .reg12        (o_d_reg[32][12]),
                .reg13        (o_d_reg[32][13]),
                .reg14        (o_d_reg[32][14]),
                .reg15        (o_d_reg[32][15]),
                .reg16        (o_d_reg[32][16]),
                .reg17        (o_d_reg[32][17]),
                .reg18        (o_d_reg[32][18]),
                .reg19        (o_d_reg[32][19]),
                .reg20        (o_d_reg[32][20]),
                .reg21        (o_d_reg[32][21]),
                .reg22        (o_d_reg[32][22]),
                .reg23        (o_d_reg[32][23]),
                .reg24        (o_d_reg[32][24]),
                .reg25        (o_d_reg[32][25]),
                .reg26        (o_d_reg[32][26]),
                .reg27        (o_d_reg[32][27]),
                .reg28        (o_d_reg[32][28]),
                .reg29        (o_d_reg[32][29]),
                .reg30        (o_d_reg[32][30]),
                .reg31        (o_d_reg[32][31]),
                .reg32        (o_d_reg[32][32]),
                .reg33        (o_d_reg[32][33]),
                .reg34        (o_d_reg[32][34]),
                .reg35        (o_d_reg[32][35]),
                .reg36        (o_d_reg[32][36]),
                .reg37        (o_d_reg[32][37]),
                .reg38        (o_d_reg[32][38]),
                .reg39        (o_d_reg[32][39]),
                .reg40        (o_d_reg[32][40]),
                .reg41        (o_d_reg[32][41]),
                .reg42        (o_d_reg[32][42]),
                .reg43        (o_d_reg[32][43]),
                .reg44        (o_d_reg[32][44]),
                .reg45        (o_d_reg[32][45]),
                .reg46        (o_d_reg[32][46]),
                .reg47        (o_d_reg[32][47]),
                .reg48        (o_d_reg[32][48]),
                .reg49        (o_d_reg[32][49]),
                .reg50        (o_d_reg[32][50]),
                .reg51        (o_d_reg[32][51]),
                .reg52        (o_d_reg[32][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf33
        (
                .din        (o_d_rowBuf[32]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[33]),
                .reg01        (o_d_reg[33][1]),
                .reg02        (o_d_reg[33][2]),
                .reg03        (o_d_reg[33][3]),
                .reg04        (o_d_reg[33][4]),
                .reg05        (o_d_reg[33][5]),
                .reg06        (o_d_reg[33][6]),
                .reg07        (o_d_reg[33][7]),
                .reg08        (o_d_reg[33][8]),
                .reg09        (o_d_reg[33][9]),
                .reg10        (o_d_reg[33][10]),
                .reg11        (o_d_reg[33][11]),
                .reg12        (o_d_reg[33][12]),
                .reg13        (o_d_reg[33][13]),
                .reg14        (o_d_reg[33][14]),
                .reg15        (o_d_reg[33][15]),
                .reg16        (o_d_reg[33][16]),
                .reg17        (o_d_reg[33][17]),
                .reg18        (o_d_reg[33][18]),
                .reg19        (o_d_reg[33][19]),
                .reg20        (o_d_reg[33][20]),
                .reg21        (o_d_reg[33][21]),
                .reg22        (o_d_reg[33][22]),
                .reg23        (o_d_reg[33][23]),
                .reg24        (o_d_reg[33][24]),
                .reg25        (o_d_reg[33][25]),
                .reg26        (o_d_reg[33][26]),
                .reg27        (o_d_reg[33][27]),
                .reg28        (o_d_reg[33][28]),
                .reg29        (o_d_reg[33][29]),
                .reg30        (o_d_reg[33][30]),
                .reg31        (o_d_reg[33][31]),
                .reg32        (o_d_reg[33][32]),
                .reg33        (o_d_reg[33][33]),
                .reg34        (o_d_reg[33][34]),
                .reg35        (o_d_reg[33][35]),
                .reg36        (o_d_reg[33][36]),
                .reg37        (o_d_reg[33][37]),
                .reg38        (o_d_reg[33][38]),
                .reg39        (o_d_reg[33][39]),
                .reg40        (o_d_reg[33][40]),
                .reg41        (o_d_reg[33][41]),
                .reg42        (o_d_reg[33][42]),
                .reg43        (o_d_reg[33][43]),
                .reg44        (o_d_reg[33][44]),
                .reg45        (o_d_reg[33][45]),
                .reg46        (o_d_reg[33][46]),
                .reg47        (o_d_reg[33][47]),
                .reg48        (o_d_reg[33][48]),
                .reg49        (o_d_reg[33][49]),
                .reg50        (o_d_reg[33][50]),
                .reg51        (o_d_reg[33][51]),
                .reg52        (o_d_reg[33][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf34
        (
                .din        (o_d_rowBuf[33]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[34]),
                .reg01        (o_d_reg[34][1]),
                .reg02        (o_d_reg[34][2]),
                .reg03        (o_d_reg[34][3]),
                .reg04        (o_d_reg[34][4]),
                .reg05        (o_d_reg[34][5]),
                .reg06        (o_d_reg[34][6]),
                .reg07        (o_d_reg[34][7]),
                .reg08        (o_d_reg[34][8]),
                .reg09        (o_d_reg[34][9]),
                .reg10        (o_d_reg[34][10]),
                .reg11        (o_d_reg[34][11]),
                .reg12        (o_d_reg[34][12]),
                .reg13        (o_d_reg[34][13]),
                .reg14        (o_d_reg[34][14]),
                .reg15        (o_d_reg[34][15]),
                .reg16        (o_d_reg[34][16]),
                .reg17        (o_d_reg[34][17]),
                .reg18        (o_d_reg[34][18]),
                .reg19        (o_d_reg[34][19]),
                .reg20        (o_d_reg[34][20]),
                .reg21        (o_d_reg[34][21]),
                .reg22        (o_d_reg[34][22]),
                .reg23        (o_d_reg[34][23]),
                .reg24        (o_d_reg[34][24]),
                .reg25        (o_d_reg[34][25]),
                .reg26        (o_d_reg[34][26]),
                .reg27        (o_d_reg[34][27]),
                .reg28        (o_d_reg[34][28]),
                .reg29        (o_d_reg[34][29]),
                .reg30        (o_d_reg[34][30]),
                .reg31        (o_d_reg[34][31]),
                .reg32        (o_d_reg[34][32]),
                .reg33        (o_d_reg[34][33]),
                .reg34        (o_d_reg[34][34]),
                .reg35        (o_d_reg[34][35]),
                .reg36        (o_d_reg[34][36]),
                .reg37        (o_d_reg[34][37]),
                .reg38        (o_d_reg[34][38]),
                .reg39        (o_d_reg[34][39]),
                .reg40        (o_d_reg[34][40]),
                .reg41        (o_d_reg[34][41]),
                .reg42        (o_d_reg[34][42]),
                .reg43        (o_d_reg[34][43]),
                .reg44        (o_d_reg[34][44]),
                .reg45        (o_d_reg[34][45]),
                .reg46        (o_d_reg[34][46]),
                .reg47        (o_d_reg[34][47]),
                .reg48        (o_d_reg[34][48]),
                .reg49        (o_d_reg[34][49]),
                .reg50        (o_d_reg[34][50]),
                .reg51        (o_d_reg[34][51]),
                .reg52        (o_d_reg[34][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf35
        (
                .din        (o_d_rowBuf[34]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[35]),
                .reg01        (o_d_reg[35][1]),
                .reg02        (o_d_reg[35][2]),
                .reg03        (o_d_reg[35][3]),
                .reg04        (o_d_reg[35][4]),
                .reg05        (o_d_reg[35][5]),
                .reg06        (o_d_reg[35][6]),
                .reg07        (o_d_reg[35][7]),
                .reg08        (o_d_reg[35][8]),
                .reg09        (o_d_reg[35][9]),
                .reg10        (o_d_reg[35][10]),
                .reg11        (o_d_reg[35][11]),
                .reg12        (o_d_reg[35][12]),
                .reg13        (o_d_reg[35][13]),
                .reg14        (o_d_reg[35][14]),
                .reg15        (o_d_reg[35][15]),
                .reg16        (o_d_reg[35][16]),
                .reg17        (o_d_reg[35][17]),
                .reg18        (o_d_reg[35][18]),
                .reg19        (o_d_reg[35][19]),
                .reg20        (o_d_reg[35][20]),
                .reg21        (o_d_reg[35][21]),
                .reg22        (o_d_reg[35][22]),
                .reg23        (o_d_reg[35][23]),
                .reg24        (o_d_reg[35][24]),
                .reg25        (o_d_reg[35][25]),
                .reg26        (o_d_reg[35][26]),
                .reg27        (o_d_reg[35][27]),
                .reg28        (o_d_reg[35][28]),
                .reg29        (o_d_reg[35][29]),
                .reg30        (o_d_reg[35][30]),
                .reg31        (o_d_reg[35][31]),
                .reg32        (o_d_reg[35][32]),
                .reg33        (o_d_reg[35][33]),
                .reg34        (o_d_reg[35][34]),
                .reg35        (o_d_reg[35][35]),
                .reg36        (o_d_reg[35][36]),
                .reg37        (o_d_reg[35][37]),
                .reg38        (o_d_reg[35][38]),
                .reg39        (o_d_reg[35][39]),
                .reg40        (o_d_reg[35][40]),
                .reg41        (o_d_reg[35][41]),
                .reg42        (o_d_reg[35][42]),
                .reg43        (o_d_reg[35][43]),
                .reg44        (o_d_reg[35][44]),
                .reg45        (o_d_reg[35][45]),
                .reg46        (o_d_reg[35][46]),
                .reg47        (o_d_reg[35][47]),
                .reg48        (o_d_reg[35][48]),
                .reg49        (o_d_reg[35][49]),
                .reg50        (o_d_reg[35][50]),
                .reg51        (o_d_reg[35][51]),
                .reg52        (o_d_reg[35][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf36
        (
                .din        (o_d_rowBuf[35]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[36]),
                .reg01        (o_d_reg[36][1]),
                .reg02        (o_d_reg[36][2]),
                .reg03        (o_d_reg[36][3]),
                .reg04        (o_d_reg[36][4]),
                .reg05        (o_d_reg[36][5]),
                .reg06        (o_d_reg[36][6]),
                .reg07        (o_d_reg[36][7]),
                .reg08        (o_d_reg[36][8]),
                .reg09        (o_d_reg[36][9]),
                .reg10        (o_d_reg[36][10]),
                .reg11        (o_d_reg[36][11]),
                .reg12        (o_d_reg[36][12]),
                .reg13        (o_d_reg[36][13]),
                .reg14        (o_d_reg[36][14]),
                .reg15        (o_d_reg[36][15]),
                .reg16        (o_d_reg[36][16]),
                .reg17        (o_d_reg[36][17]),
                .reg18        (o_d_reg[36][18]),
                .reg19        (o_d_reg[36][19]),
                .reg20        (o_d_reg[36][20]),
                .reg21        (o_d_reg[36][21]),
                .reg22        (o_d_reg[36][22]),
                .reg23        (o_d_reg[36][23]),
                .reg24        (o_d_reg[36][24]),
                .reg25        (o_d_reg[36][25]),
                .reg26        (o_d_reg[36][26]),
                .reg27        (o_d_reg[36][27]),
                .reg28        (o_d_reg[36][28]),
                .reg29        (o_d_reg[36][29]),
                .reg30        (o_d_reg[36][30]),
                .reg31        (o_d_reg[36][31]),
                .reg32        (o_d_reg[36][32]),
                .reg33        (o_d_reg[36][33]),
                .reg34        (o_d_reg[36][34]),
                .reg35        (o_d_reg[36][35]),
                .reg36        (o_d_reg[36][36]),
                .reg37        (o_d_reg[36][37]),
                .reg38        (o_d_reg[36][38]),
                .reg39        (o_d_reg[36][39]),
                .reg40        (o_d_reg[36][40]),
                .reg41        (o_d_reg[36][41]),
                .reg42        (o_d_reg[36][42]),
                .reg43        (o_d_reg[36][43]),
                .reg44        (o_d_reg[36][44]),
                .reg45        (o_d_reg[36][45]),
                .reg46        (o_d_reg[36][46]),
                .reg47        (o_d_reg[36][47]),
                .reg48        (o_d_reg[36][48]),
                .reg49        (o_d_reg[36][49]),
                .reg50        (o_d_reg[36][50]),
                .reg51        (o_d_reg[36][51]),
                .reg52        (o_d_reg[36][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf37
        (
                .din        (o_d_rowBuf[36]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[37]),
                .reg01        (o_d_reg[37][1]),
                .reg02        (o_d_reg[37][2]),
                .reg03        (o_d_reg[37][3]),
                .reg04        (o_d_reg[37][4]),
                .reg05        (o_d_reg[37][5]),
                .reg06        (o_d_reg[37][6]),
                .reg07        (o_d_reg[37][7]),
                .reg08        (o_d_reg[37][8]),
                .reg09        (o_d_reg[37][9]),
                .reg10        (o_d_reg[37][10]),
                .reg11        (o_d_reg[37][11]),
                .reg12        (o_d_reg[37][12]),
                .reg13        (o_d_reg[37][13]),
                .reg14        (o_d_reg[37][14]),
                .reg15        (o_d_reg[37][15]),
                .reg16        (o_d_reg[37][16]),
                .reg17        (o_d_reg[37][17]),
                .reg18        (o_d_reg[37][18]),
                .reg19        (o_d_reg[37][19]),
                .reg20        (o_d_reg[37][20]),
                .reg21        (o_d_reg[37][21]),
                .reg22        (o_d_reg[37][22]),
                .reg23        (o_d_reg[37][23]),
                .reg24        (o_d_reg[37][24]),
                .reg25        (o_d_reg[37][25]),
                .reg26        (o_d_reg[37][26]),
                .reg27        (o_d_reg[37][27]),
                .reg28        (o_d_reg[37][28]),
                .reg29        (o_d_reg[37][29]),
                .reg30        (o_d_reg[37][30]),
                .reg31        (o_d_reg[37][31]),
                .reg32        (o_d_reg[37][32]),
                .reg33        (o_d_reg[37][33]),
                .reg34        (o_d_reg[37][34]),
                .reg35        (o_d_reg[37][35]),
                .reg36        (o_d_reg[37][36]),
                .reg37        (o_d_reg[37][37]),
                .reg38        (o_d_reg[37][38]),
                .reg39        (o_d_reg[37][39]),
                .reg40        (o_d_reg[37][40]),
                .reg41        (o_d_reg[37][41]),
                .reg42        (o_d_reg[37][42]),
                .reg43        (o_d_reg[37][43]),
                .reg44        (o_d_reg[37][44]),
                .reg45        (o_d_reg[37][45]),
                .reg46        (o_d_reg[37][46]),
                .reg47        (o_d_reg[37][47]),
                .reg48        (o_d_reg[37][48]),
                .reg49        (o_d_reg[37][49]),
                .reg50        (o_d_reg[37][50]),
                .reg51        (o_d_reg[37][51]),
                .reg52        (o_d_reg[37][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf38
        (
                .din        (o_d_rowBuf[37]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[38]),
                .reg01        (o_d_reg[38][1]),
                .reg02        (o_d_reg[38][2]),
                .reg03        (o_d_reg[38][3]),
                .reg04        (o_d_reg[38][4]),
                .reg05        (o_d_reg[38][5]),
                .reg06        (o_d_reg[38][6]),
                .reg07        (o_d_reg[38][7]),
                .reg08        (o_d_reg[38][8]),
                .reg09        (o_d_reg[38][9]),
                .reg10        (o_d_reg[38][10]),
                .reg11        (o_d_reg[38][11]),
                .reg12        (o_d_reg[38][12]),
                .reg13        (o_d_reg[38][13]),
                .reg14        (o_d_reg[38][14]),
                .reg15        (o_d_reg[38][15]),
                .reg16        (o_d_reg[38][16]),
                .reg17        (o_d_reg[38][17]),
                .reg18        (o_d_reg[38][18]),
                .reg19        (o_d_reg[38][19]),
                .reg20        (o_d_reg[38][20]),
                .reg21        (o_d_reg[38][21]),
                .reg22        (o_d_reg[38][22]),
                .reg23        (o_d_reg[38][23]),
                .reg24        (o_d_reg[38][24]),
                .reg25        (o_d_reg[38][25]),
                .reg26        (o_d_reg[38][26]),
                .reg27        (o_d_reg[38][27]),
                .reg28        (o_d_reg[38][28]),
                .reg29        (o_d_reg[38][29]),
                .reg30        (o_d_reg[38][30]),
                .reg31        (o_d_reg[38][31]),
                .reg32        (o_d_reg[38][32]),
                .reg33        (o_d_reg[38][33]),
                .reg34        (o_d_reg[38][34]),
                .reg35        (o_d_reg[38][35]),
                .reg36        (o_d_reg[38][36]),
                .reg37        (o_d_reg[38][37]),
                .reg38        (o_d_reg[38][38]),
                .reg39        (o_d_reg[38][39]),
                .reg40        (o_d_reg[38][40]),
                .reg41        (o_d_reg[38][41]),
                .reg42        (o_d_reg[38][42]),
                .reg43        (o_d_reg[38][43]),
                .reg44        (o_d_reg[38][44]),
                .reg45        (o_d_reg[38][45]),
                .reg46        (o_d_reg[38][46]),
                .reg47        (o_d_reg[38][47]),
                .reg48        (o_d_reg[38][48]),
                .reg49        (o_d_reg[38][49]),
                .reg50        (o_d_reg[38][50]),
                .reg51        (o_d_reg[38][51]),
                .reg52        (o_d_reg[38][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf39
        (
                .din        (o_d_rowBuf[38]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[39]),
                .reg01        (o_d_reg[39][1]),
                .reg02        (o_d_reg[39][2]),
                .reg03        (o_d_reg[39][3]),
                .reg04        (o_d_reg[39][4]),
                .reg05        (o_d_reg[39][5]),
                .reg06        (o_d_reg[39][6]),
                .reg07        (o_d_reg[39][7]),
                .reg08        (o_d_reg[39][8]),
                .reg09        (o_d_reg[39][9]),
                .reg10        (o_d_reg[39][10]),
                .reg11        (o_d_reg[39][11]),
                .reg12        (o_d_reg[39][12]),
                .reg13        (o_d_reg[39][13]),
                .reg14        (o_d_reg[39][14]),
                .reg15        (o_d_reg[39][15]),
                .reg16        (o_d_reg[39][16]),
                .reg17        (o_d_reg[39][17]),
                .reg18        (o_d_reg[39][18]),
                .reg19        (o_d_reg[39][19]),
                .reg20        (o_d_reg[39][20]),
                .reg21        (o_d_reg[39][21]),
                .reg22        (o_d_reg[39][22]),
                .reg23        (o_d_reg[39][23]),
                .reg24        (o_d_reg[39][24]),
                .reg25        (o_d_reg[39][25]),
                .reg26        (o_d_reg[39][26]),
                .reg27        (o_d_reg[39][27]),
                .reg28        (o_d_reg[39][28]),
                .reg29        (o_d_reg[39][29]),
                .reg30        (o_d_reg[39][30]),
                .reg31        (o_d_reg[39][31]),
                .reg32        (o_d_reg[39][32]),
                .reg33        (o_d_reg[39][33]),
                .reg34        (o_d_reg[39][34]),
                .reg35        (o_d_reg[39][35]),
                .reg36        (o_d_reg[39][36]),
                .reg37        (o_d_reg[39][37]),
                .reg38        (o_d_reg[39][38]),
                .reg39        (o_d_reg[39][39]),
                .reg40        (o_d_reg[39][40]),
                .reg41        (o_d_reg[39][41]),
                .reg42        (o_d_reg[39][42]),
                .reg43        (o_d_reg[39][43]),
                .reg44        (o_d_reg[39][44]),
                .reg45        (o_d_reg[39][45]),
                .reg46        (o_d_reg[39][46]),
                .reg47        (o_d_reg[39][47]),
                .reg48        (o_d_reg[39][48]),
                .reg49        (o_d_reg[39][49]),
                .reg50        (o_d_reg[39][50]),
                .reg51        (o_d_reg[39][51]),
                .reg52        (o_d_reg[39][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf40
        (
                .din        (o_d_rowBuf[39]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[40]),
                .reg01        (o_d_reg[40][1]),
                .reg02        (o_d_reg[40][2]),
                .reg03        (o_d_reg[40][3]),
                .reg04        (o_d_reg[40][4]),
                .reg05        (o_d_reg[40][5]),
                .reg06        (o_d_reg[40][6]),
                .reg07        (o_d_reg[40][7]),
                .reg08        (o_d_reg[40][8]),
                .reg09        (o_d_reg[40][9]),
                .reg10        (o_d_reg[40][10]),
                .reg11        (o_d_reg[40][11]),
                .reg12        (o_d_reg[40][12]),
                .reg13        (o_d_reg[40][13]),
                .reg14        (o_d_reg[40][14]),
                .reg15        (o_d_reg[40][15]),
                .reg16        (o_d_reg[40][16]),
                .reg17        (o_d_reg[40][17]),
                .reg18        (o_d_reg[40][18]),
                .reg19        (o_d_reg[40][19]),
                .reg20        (o_d_reg[40][20]),
                .reg21        (o_d_reg[40][21]),
                .reg22        (o_d_reg[40][22]),
                .reg23        (o_d_reg[40][23]),
                .reg24        (o_d_reg[40][24]),
                .reg25        (o_d_reg[40][25]),
                .reg26        (o_d_reg[40][26]),
                .reg27        (o_d_reg[40][27]),
                .reg28        (o_d_reg[40][28]),
                .reg29        (o_d_reg[40][29]),
                .reg30        (o_d_reg[40][30]),
                .reg31        (o_d_reg[40][31]),
                .reg32        (o_d_reg[40][32]),
                .reg33        (o_d_reg[40][33]),
                .reg34        (o_d_reg[40][34]),
                .reg35        (o_d_reg[40][35]),
                .reg36        (o_d_reg[40][36]),
                .reg37        (o_d_reg[40][37]),
                .reg38        (o_d_reg[40][38]),
                .reg39        (o_d_reg[40][39]),
                .reg40        (o_d_reg[40][40]),
                .reg41        (o_d_reg[40][41]),
                .reg42        (o_d_reg[40][42]),
                .reg43        (o_d_reg[40][43]),
                .reg44        (o_d_reg[40][44]),
                .reg45        (o_d_reg[40][45]),
                .reg46        (o_d_reg[40][46]),
                .reg47        (o_d_reg[40][47]),
                .reg48        (o_d_reg[40][48]),
                .reg49        (o_d_reg[40][49]),
                .reg50        (o_d_reg[40][50]),
                .reg51        (o_d_reg[40][51]),
                .reg52        (o_d_reg[40][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf41
        (
                .din        (o_d_rowBuf[40]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[41]),
                .reg01        (o_d_reg[41][1]),
                .reg02        (o_d_reg[41][2]),
                .reg03        (o_d_reg[41][3]),
                .reg04        (o_d_reg[41][4]),
                .reg05        (o_d_reg[41][5]),
                .reg06        (o_d_reg[41][6]),
                .reg07        (o_d_reg[41][7]),
                .reg08        (o_d_reg[41][8]),
                .reg09        (o_d_reg[41][9]),
                .reg10        (o_d_reg[41][10]),
                .reg11        (o_d_reg[41][11]),
                .reg12        (o_d_reg[41][12]),
                .reg13        (o_d_reg[41][13]),
                .reg14        (o_d_reg[41][14]),
                .reg15        (o_d_reg[41][15]),
                .reg16        (o_d_reg[41][16]),
                .reg17        (o_d_reg[41][17]),
                .reg18        (o_d_reg[41][18]),
                .reg19        (o_d_reg[41][19]),
                .reg20        (o_d_reg[41][20]),
                .reg21        (o_d_reg[41][21]),
                .reg22        (o_d_reg[41][22]),
                .reg23        (o_d_reg[41][23]),
                .reg24        (o_d_reg[41][24]),
                .reg25        (o_d_reg[41][25]),
                .reg26        (o_d_reg[41][26]),
                .reg27        (o_d_reg[41][27]),
                .reg28        (o_d_reg[41][28]),
                .reg29        (o_d_reg[41][29]),
                .reg30        (o_d_reg[41][30]),
                .reg31        (o_d_reg[41][31]),
                .reg32        (o_d_reg[41][32]),
                .reg33        (o_d_reg[41][33]),
                .reg34        (o_d_reg[41][34]),
                .reg35        (o_d_reg[41][35]),
                .reg36        (o_d_reg[41][36]),
                .reg37        (o_d_reg[41][37]),
                .reg38        (o_d_reg[41][38]),
                .reg39        (o_d_reg[41][39]),
                .reg40        (o_d_reg[41][40]),
                .reg41        (o_d_reg[41][41]),
                .reg42        (o_d_reg[41][42]),
                .reg43        (o_d_reg[41][43]),
                .reg44        (o_d_reg[41][44]),
                .reg45        (o_d_reg[41][45]),
                .reg46        (o_d_reg[41][46]),
                .reg47        (o_d_reg[41][47]),
                .reg48        (o_d_reg[41][48]),
                .reg49        (o_d_reg[41][49]),
                .reg50        (o_d_reg[41][50]),
                .reg51        (o_d_reg[41][51]),
                .reg52        (o_d_reg[41][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf42
        (
                .din        (o_d_rowBuf[41]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[42]),
                .reg01        (o_d_reg[42][1]),
                .reg02        (o_d_reg[42][2]),
                .reg03        (o_d_reg[42][3]),
                .reg04        (o_d_reg[42][4]),
                .reg05        (o_d_reg[42][5]),
                .reg06        (o_d_reg[42][6]),
                .reg07        (o_d_reg[42][7]),
                .reg08        (o_d_reg[42][8]),
                .reg09        (o_d_reg[42][9]),
                .reg10        (o_d_reg[42][10]),
                .reg11        (o_d_reg[42][11]),
                .reg12        (o_d_reg[42][12]),
                .reg13        (o_d_reg[42][13]),
                .reg14        (o_d_reg[42][14]),
                .reg15        (o_d_reg[42][15]),
                .reg16        (o_d_reg[42][16]),
                .reg17        (o_d_reg[42][17]),
                .reg18        (o_d_reg[42][18]),
                .reg19        (o_d_reg[42][19]),
                .reg20        (o_d_reg[42][20]),
                .reg21        (o_d_reg[42][21]),
                .reg22        (o_d_reg[42][22]),
                .reg23        (o_d_reg[42][23]),
                .reg24        (o_d_reg[42][24]),
                .reg25        (o_d_reg[42][25]),
                .reg26        (o_d_reg[42][26]),
                .reg27        (o_d_reg[42][27]),
                .reg28        (o_d_reg[42][28]),
                .reg29        (o_d_reg[42][29]),
                .reg30        (o_d_reg[42][30]),
                .reg31        (o_d_reg[42][31]),
                .reg32        (o_d_reg[42][32]),
                .reg33        (o_d_reg[42][33]),
                .reg34        (o_d_reg[42][34]),
                .reg35        (o_d_reg[42][35]),
                .reg36        (o_d_reg[42][36]),
                .reg37        (o_d_reg[42][37]),
                .reg38        (o_d_reg[42][38]),
                .reg39        (o_d_reg[42][39]),
                .reg40        (o_d_reg[42][40]),
                .reg41        (o_d_reg[42][41]),
                .reg42        (o_d_reg[42][42]),
                .reg43        (o_d_reg[42][43]),
                .reg44        (o_d_reg[42][44]),
                .reg45        (o_d_reg[42][45]),
                .reg46        (o_d_reg[42][46]),
                .reg47        (o_d_reg[42][47]),
                .reg48        (o_d_reg[42][48]),
                .reg49        (o_d_reg[42][49]),
                .reg50        (o_d_reg[42][50]),
                .reg51        (o_d_reg[42][51]),
                .reg52        (o_d_reg[42][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf43
        (
                .din        (o_d_rowBuf[42]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[43]),
                .reg01        (o_d_reg[43][1]),
                .reg02        (o_d_reg[43][2]),
                .reg03        (o_d_reg[43][3]),
                .reg04        (o_d_reg[43][4]),
                .reg05        (o_d_reg[43][5]),
                .reg06        (o_d_reg[43][6]),
                .reg07        (o_d_reg[43][7]),
                .reg08        (o_d_reg[43][8]),
                .reg09        (o_d_reg[43][9]),
                .reg10        (o_d_reg[43][10]),
                .reg11        (o_d_reg[43][11]),
                .reg12        (o_d_reg[43][12]),
                .reg13        (o_d_reg[43][13]),
                .reg14        (o_d_reg[43][14]),
                .reg15        (o_d_reg[43][15]),
                .reg16        (o_d_reg[43][16]),
                .reg17        (o_d_reg[43][17]),
                .reg18        (o_d_reg[43][18]),
                .reg19        (o_d_reg[43][19]),
                .reg20        (o_d_reg[43][20]),
                .reg21        (o_d_reg[43][21]),
                .reg22        (o_d_reg[43][22]),
                .reg23        (o_d_reg[43][23]),
                .reg24        (o_d_reg[43][24]),
                .reg25        (o_d_reg[43][25]),
                .reg26        (o_d_reg[43][26]),
                .reg27        (o_d_reg[43][27]),
                .reg28        (o_d_reg[43][28]),
                .reg29        (o_d_reg[43][29]),
                .reg30        (o_d_reg[43][30]),
                .reg31        (o_d_reg[43][31]),
                .reg32        (o_d_reg[43][32]),
                .reg33        (o_d_reg[43][33]),
                .reg34        (o_d_reg[43][34]),
                .reg35        (o_d_reg[43][35]),
                .reg36        (o_d_reg[43][36]),
                .reg37        (o_d_reg[43][37]),
                .reg38        (o_d_reg[43][38]),
                .reg39        (o_d_reg[43][39]),
                .reg40        (o_d_reg[43][40]),
                .reg41        (o_d_reg[43][41]),
                .reg42        (o_d_reg[43][42]),
                .reg43        (o_d_reg[43][43]),
                .reg44        (o_d_reg[43][44]),
                .reg45        (o_d_reg[43][45]),
                .reg46        (o_d_reg[43][46]),
                .reg47        (o_d_reg[43][47]),
                .reg48        (o_d_reg[43][48]),
                .reg49        (o_d_reg[43][49]),
                .reg50        (o_d_reg[43][50]),
                .reg51        (o_d_reg[43][51]),
                .reg52        (o_d_reg[43][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf44
        (
                .din        (o_d_rowBuf[43]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[44]),
                .reg01        (o_d_reg[44][1]),
                .reg02        (o_d_reg[44][2]),
                .reg03        (o_d_reg[44][3]),
                .reg04        (o_d_reg[44][4]),
                .reg05        (o_d_reg[44][5]),
                .reg06        (o_d_reg[44][6]),
                .reg07        (o_d_reg[44][7]),
                .reg08        (o_d_reg[44][8]),
                .reg09        (o_d_reg[44][9]),
                .reg10        (o_d_reg[44][10]),
                .reg11        (o_d_reg[44][11]),
                .reg12        (o_d_reg[44][12]),
                .reg13        (o_d_reg[44][13]),
                .reg14        (o_d_reg[44][14]),
                .reg15        (o_d_reg[44][15]),
                .reg16        (o_d_reg[44][16]),
                .reg17        (o_d_reg[44][17]),
                .reg18        (o_d_reg[44][18]),
                .reg19        (o_d_reg[44][19]),
                .reg20        (o_d_reg[44][20]),
                .reg21        (o_d_reg[44][21]),
                .reg22        (o_d_reg[44][22]),
                .reg23        (o_d_reg[44][23]),
                .reg24        (o_d_reg[44][24]),
                .reg25        (o_d_reg[44][25]),
                .reg26        (o_d_reg[44][26]),
                .reg27        (o_d_reg[44][27]),
                .reg28        (o_d_reg[44][28]),
                .reg29        (o_d_reg[44][29]),
                .reg30        (o_d_reg[44][30]),
                .reg31        (o_d_reg[44][31]),
                .reg32        (o_d_reg[44][32]),
                .reg33        (o_d_reg[44][33]),
                .reg34        (o_d_reg[44][34]),
                .reg35        (o_d_reg[44][35]),
                .reg36        (o_d_reg[44][36]),
                .reg37        (o_d_reg[44][37]),
                .reg38        (o_d_reg[44][38]),
                .reg39        (o_d_reg[44][39]),
                .reg40        (o_d_reg[44][40]),
                .reg41        (o_d_reg[44][41]),
                .reg42        (o_d_reg[44][42]),
                .reg43        (o_d_reg[44][43]),
                .reg44        (o_d_reg[44][44]),
                .reg45        (o_d_reg[44][45]),
                .reg46        (o_d_reg[44][46]),
                .reg47        (o_d_reg[44][47]),
                .reg48        (o_d_reg[44][48]),
                .reg49        (o_d_reg[44][49]),
                .reg50        (o_d_reg[44][50]),
                .reg51        (o_d_reg[44][51]),
                .reg52        (o_d_reg[44][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf45
        (
                .din        (o_d_rowBuf[44]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[45]),
                .reg01        (o_d_reg[45][1]),
                .reg02        (o_d_reg[45][2]),
                .reg03        (o_d_reg[45][3]),
                .reg04        (o_d_reg[45][4]),
                .reg05        (o_d_reg[45][5]),
                .reg06        (o_d_reg[45][6]),
                .reg07        (o_d_reg[45][7]),
                .reg08        (o_d_reg[45][8]),
                .reg09        (o_d_reg[45][9]),
                .reg10        (o_d_reg[45][10]),
                .reg11        (o_d_reg[45][11]),
                .reg12        (o_d_reg[45][12]),
                .reg13        (o_d_reg[45][13]),
                .reg14        (o_d_reg[45][14]),
                .reg15        (o_d_reg[45][15]),
                .reg16        (o_d_reg[45][16]),
                .reg17        (o_d_reg[45][17]),
                .reg18        (o_d_reg[45][18]),
                .reg19        (o_d_reg[45][19]),
                .reg20        (o_d_reg[45][20]),
                .reg21        (o_d_reg[45][21]),
                .reg22        (o_d_reg[45][22]),
                .reg23        (o_d_reg[45][23]),
                .reg24        (o_d_reg[45][24]),
                .reg25        (o_d_reg[45][25]),
                .reg26        (o_d_reg[45][26]),
                .reg27        (o_d_reg[45][27]),
                .reg28        (o_d_reg[45][28]),
                .reg29        (o_d_reg[45][29]),
                .reg30        (o_d_reg[45][30]),
                .reg31        (o_d_reg[45][31]),
                .reg32        (o_d_reg[45][32]),
                .reg33        (o_d_reg[45][33]),
                .reg34        (o_d_reg[45][34]),
                .reg35        (o_d_reg[45][35]),
                .reg36        (o_d_reg[45][36]),
                .reg37        (o_d_reg[45][37]),
                .reg38        (o_d_reg[45][38]),
                .reg39        (o_d_reg[45][39]),
                .reg40        (o_d_reg[45][40]),
                .reg41        (o_d_reg[45][41]),
                .reg42        (o_d_reg[45][42]),
                .reg43        (o_d_reg[45][43]),
                .reg44        (o_d_reg[45][44]),
                .reg45        (o_d_reg[45][45]),
                .reg46        (o_d_reg[45][46]),
                .reg47        (o_d_reg[45][47]),
                .reg48        (o_d_reg[45][48]),
                .reg49        (o_d_reg[45][49]),
                .reg50        (o_d_reg[45][50]),
                .reg51        (o_d_reg[45][51]),
                .reg52        (o_d_reg[45][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf46
        (
                .din        (o_d_rowBuf[45]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[46]),
                .reg01        (o_d_reg[46][1]),
                .reg02        (o_d_reg[46][2]),
                .reg03        (o_d_reg[46][3]),
                .reg04        (o_d_reg[46][4]),
                .reg05        (o_d_reg[46][5]),
                .reg06        (o_d_reg[46][6]),
                .reg07        (o_d_reg[46][7]),
                .reg08        (o_d_reg[46][8]),
                .reg09        (o_d_reg[46][9]),
                .reg10        (o_d_reg[46][10]),
                .reg11        (o_d_reg[46][11]),
                .reg12        (o_d_reg[46][12]),
                .reg13        (o_d_reg[46][13]),
                .reg14        (o_d_reg[46][14]),
                .reg15        (o_d_reg[46][15]),
                .reg16        (o_d_reg[46][16]),
                .reg17        (o_d_reg[46][17]),
                .reg18        (o_d_reg[46][18]),
                .reg19        (o_d_reg[46][19]),
                .reg20        (o_d_reg[46][20]),
                .reg21        (o_d_reg[46][21]),
                .reg22        (o_d_reg[46][22]),
                .reg23        (o_d_reg[46][23]),
                .reg24        (o_d_reg[46][24]),
                .reg25        (o_d_reg[46][25]),
                .reg26        (o_d_reg[46][26]),
                .reg27        (o_d_reg[46][27]),
                .reg28        (o_d_reg[46][28]),
                .reg29        (o_d_reg[46][29]),
                .reg30        (o_d_reg[46][30]),
                .reg31        (o_d_reg[46][31]),
                .reg32        (o_d_reg[46][32]),
                .reg33        (o_d_reg[46][33]),
                .reg34        (o_d_reg[46][34]),
                .reg35        (o_d_reg[46][35]),
                .reg36        (o_d_reg[46][36]),
                .reg37        (o_d_reg[46][37]),
                .reg38        (o_d_reg[46][38]),
                .reg39        (o_d_reg[46][39]),
                .reg40        (o_d_reg[46][40]),
                .reg41        (o_d_reg[46][41]),
                .reg42        (o_d_reg[46][42]),
                .reg43        (o_d_reg[46][43]),
                .reg44        (o_d_reg[46][44]),
                .reg45        (o_d_reg[46][45]),
                .reg46        (o_d_reg[46][46]),
                .reg47        (o_d_reg[46][47]),
                .reg48        (o_d_reg[46][48]),
                .reg49        (o_d_reg[46][49]),
                .reg50        (o_d_reg[46][50]),
                .reg51        (o_d_reg[46][51]),
                .reg52        (o_d_reg[46][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf47
        (
                .din        (o_d_rowBuf[46]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[47]),
                .reg01        (o_d_reg[47][1]),
                .reg02        (o_d_reg[47][2]),
                .reg03        (o_d_reg[47][3]),
                .reg04        (o_d_reg[47][4]),
                .reg05        (o_d_reg[47][5]),
                .reg06        (o_d_reg[47][6]),
                .reg07        (o_d_reg[47][7]),
                .reg08        (o_d_reg[47][8]),
                .reg09        (o_d_reg[47][9]),
                .reg10        (o_d_reg[47][10]),
                .reg11        (o_d_reg[47][11]),
                .reg12        (o_d_reg[47][12]),
                .reg13        (o_d_reg[47][13]),
                .reg14        (o_d_reg[47][14]),
                .reg15        (o_d_reg[47][15]),
                .reg16        (o_d_reg[47][16]),
                .reg17        (o_d_reg[47][17]),
                .reg18        (o_d_reg[47][18]),
                .reg19        (o_d_reg[47][19]),
                .reg20        (o_d_reg[47][20]),
                .reg21        (o_d_reg[47][21]),
                .reg22        (o_d_reg[47][22]),
                .reg23        (o_d_reg[47][23]),
                .reg24        (o_d_reg[47][24]),
                .reg25        (o_d_reg[47][25]),
                .reg26        (o_d_reg[47][26]),
                .reg27        (o_d_reg[47][27]),
                .reg28        (o_d_reg[47][28]),
                .reg29        (o_d_reg[47][29]),
                .reg30        (o_d_reg[47][30]),
                .reg31        (o_d_reg[47][31]),
                .reg32        (o_d_reg[47][32]),
                .reg33        (o_d_reg[47][33]),
                .reg34        (o_d_reg[47][34]),
                .reg35        (o_d_reg[47][35]),
                .reg36        (o_d_reg[47][36]),
                .reg37        (o_d_reg[47][37]),
                .reg38        (o_d_reg[47][38]),
                .reg39        (o_d_reg[47][39]),
                .reg40        (o_d_reg[47][40]),
                .reg41        (o_d_reg[47][41]),
                .reg42        (o_d_reg[47][42]),
                .reg43        (o_d_reg[47][43]),
                .reg44        (o_d_reg[47][44]),
                .reg45        (o_d_reg[47][45]),
                .reg46        (o_d_reg[47][46]),
                .reg47        (o_d_reg[47][47]),
                .reg48        (o_d_reg[47][48]),
                .reg49        (o_d_reg[47][49]),
                .reg50        (o_d_reg[47][50]),
                .reg51        (o_d_reg[47][51]),
                .reg52        (o_d_reg[47][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf48
        (
                .din        (o_d_rowBuf[47]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[48]),
                .reg01        (o_d_reg[48][1]),
                .reg02        (o_d_reg[48][2]),
                .reg03        (o_d_reg[48][3]),
                .reg04        (o_d_reg[48][4]),
                .reg05        (o_d_reg[48][5]),
                .reg06        (o_d_reg[48][6]),
                .reg07        (o_d_reg[48][7]),
                .reg08        (o_d_reg[48][8]),
                .reg09        (o_d_reg[48][9]),
                .reg10        (o_d_reg[48][10]),
                .reg11        (o_d_reg[48][11]),
                .reg12        (o_d_reg[48][12]),
                .reg13        (o_d_reg[48][13]),
                .reg14        (o_d_reg[48][14]),
                .reg15        (o_d_reg[48][15]),
                .reg16        (o_d_reg[48][16]),
                .reg17        (o_d_reg[48][17]),
                .reg18        (o_d_reg[48][18]),
                .reg19        (o_d_reg[48][19]),
                .reg20        (o_d_reg[48][20]),
                .reg21        (o_d_reg[48][21]),
                .reg22        (o_d_reg[48][22]),
                .reg23        (o_d_reg[48][23]),
                .reg24        (o_d_reg[48][24]),
                .reg25        (o_d_reg[48][25]),
                .reg26        (o_d_reg[48][26]),
                .reg27        (o_d_reg[48][27]),
                .reg28        (o_d_reg[48][28]),
                .reg29        (o_d_reg[48][29]),
                .reg30        (o_d_reg[48][30]),
                .reg31        (o_d_reg[48][31]),
                .reg32        (o_d_reg[48][32]),
                .reg33        (o_d_reg[48][33]),
                .reg34        (o_d_reg[48][34]),
                .reg35        (o_d_reg[48][35]),
                .reg36        (o_d_reg[48][36]),
                .reg37        (o_d_reg[48][37]),
                .reg38        (o_d_reg[48][38]),
                .reg39        (o_d_reg[48][39]),
                .reg40        (o_d_reg[48][40]),
                .reg41        (o_d_reg[48][41]),
                .reg42        (o_d_reg[48][42]),
                .reg43        (o_d_reg[48][43]),
                .reg44        (o_d_reg[48][44]),
                .reg45        (o_d_reg[48][45]),
                .reg46        (o_d_reg[48][46]),
                .reg47        (o_d_reg[48][47]),
                .reg48        (o_d_reg[48][48]),
                .reg49        (o_d_reg[48][49]),
                .reg50        (o_d_reg[48][50]),
                .reg51        (o_d_reg[48][51]),
                .reg52        (o_d_reg[48][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf49
        (
                .din        (o_d_rowBuf[48]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[49]),
                .reg01        (o_d_reg[49][1]),
                .reg02        (o_d_reg[49][2]),
                .reg03        (o_d_reg[49][3]),
                .reg04        (o_d_reg[49][4]),
                .reg05        (o_d_reg[49][5]),
                .reg06        (o_d_reg[49][6]),
                .reg07        (o_d_reg[49][7]),
                .reg08        (o_d_reg[49][8]),
                .reg09        (o_d_reg[49][9]),
                .reg10        (o_d_reg[49][10]),
                .reg11        (o_d_reg[49][11]),
                .reg12        (o_d_reg[49][12]),
                .reg13        (o_d_reg[49][13]),
                .reg14        (o_d_reg[49][14]),
                .reg15        (o_d_reg[49][15]),
                .reg16        (o_d_reg[49][16]),
                .reg17        (o_d_reg[49][17]),
                .reg18        (o_d_reg[49][18]),
                .reg19        (o_d_reg[49][19]),
                .reg20        (o_d_reg[49][20]),
                .reg21        (o_d_reg[49][21]),
                .reg22        (o_d_reg[49][22]),
                .reg23        (o_d_reg[49][23]),
                .reg24        (o_d_reg[49][24]),
                .reg25        (o_d_reg[49][25]),
                .reg26        (o_d_reg[49][26]),
                .reg27        (o_d_reg[49][27]),
                .reg28        (o_d_reg[49][28]),
                .reg29        (o_d_reg[49][29]),
                .reg30        (o_d_reg[49][30]),
                .reg31        (o_d_reg[49][31]),
                .reg32        (o_d_reg[49][32]),
                .reg33        (o_d_reg[49][33]),
                .reg34        (o_d_reg[49][34]),
                .reg35        (o_d_reg[49][35]),
                .reg36        (o_d_reg[49][36]),
                .reg37        (o_d_reg[49][37]),
                .reg38        (o_d_reg[49][38]),
                .reg39        (o_d_reg[49][39]),
                .reg40        (o_d_reg[49][40]),
                .reg41        (o_d_reg[49][41]),
                .reg42        (o_d_reg[49][42]),
                .reg43        (o_d_reg[49][43]),
                .reg44        (o_d_reg[49][44]),
                .reg45        (o_d_reg[49][45]),
                .reg46        (o_d_reg[49][46]),
                .reg47        (o_d_reg[49][47]),
                .reg48        (o_d_reg[49][48]),
                .reg49        (o_d_reg[49][49]),
                .reg50        (o_d_reg[49][50]),
                .reg51        (o_d_reg[49][51]),
                .reg52        (o_d_reg[49][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf50
        (
                .din        (o_d_rowBuf[49]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[50]),
                .reg01        (o_d_reg[50][1]),
                .reg02        (o_d_reg[50][2]),
                .reg03        (o_d_reg[50][3]),
                .reg04        (o_d_reg[50][4]),
                .reg05        (o_d_reg[50][5]),
                .reg06        (o_d_reg[50][6]),
                .reg07        (o_d_reg[50][7]),
                .reg08        (o_d_reg[50][8]),
                .reg09        (o_d_reg[50][9]),
                .reg10        (o_d_reg[50][10]),
                .reg11        (o_d_reg[50][11]),
                .reg12        (o_d_reg[50][12]),
                .reg13        (o_d_reg[50][13]),
                .reg14        (o_d_reg[50][14]),
                .reg15        (o_d_reg[50][15]),
                .reg16        (o_d_reg[50][16]),
                .reg17        (o_d_reg[50][17]),
                .reg18        (o_d_reg[50][18]),
                .reg19        (o_d_reg[50][19]),
                .reg20        (o_d_reg[50][20]),
                .reg21        (o_d_reg[50][21]),
                .reg22        (o_d_reg[50][22]),
                .reg23        (o_d_reg[50][23]),
                .reg24        (o_d_reg[50][24]),
                .reg25        (o_d_reg[50][25]),
                .reg26        (o_d_reg[50][26]),
                .reg27        (o_d_reg[50][27]),
                .reg28        (o_d_reg[50][28]),
                .reg29        (o_d_reg[50][29]),
                .reg30        (o_d_reg[50][30]),
                .reg31        (o_d_reg[50][31]),
                .reg32        (o_d_reg[50][32]),
                .reg33        (o_d_reg[50][33]),
                .reg34        (o_d_reg[50][34]),
                .reg35        (o_d_reg[50][35]),
                .reg36        (o_d_reg[50][36]),
                .reg37        (o_d_reg[50][37]),
                .reg38        (o_d_reg[50][38]),
                .reg39        (o_d_reg[50][39]),
                .reg40        (o_d_reg[50][40]),
                .reg41        (o_d_reg[50][41]),
                .reg42        (o_d_reg[50][42]),
                .reg43        (o_d_reg[50][43]),
                .reg44        (o_d_reg[50][44]),
                .reg45        (o_d_reg[50][45]),
                .reg46        (o_d_reg[50][46]),
                .reg47        (o_d_reg[50][47]),
                .reg48        (o_d_reg[50][48]),
                .reg49        (o_d_reg[50][49]),
                .reg50        (o_d_reg[50][50]),
                .reg51        (o_d_reg[50][51]),
                .reg52        (o_d_reg[50][52])
        );
        rowBuf #(.IMAGE_WIDTH (IMAGE_WIDTH))	rowBuf51
        (
                .din        (o_d_rowBuf[50]),
                .clk        (clk),
                .rst        (rst),
                .dout        (o_d_rowBuf[51]),
                .reg01        (o_d_reg[51][1]),
                .reg02        (o_d_reg[51][2]),
                .reg03        (o_d_reg[51][3]),
                .reg04        (o_d_reg[51][4]),
                .reg05        (o_d_reg[51][5]),
                .reg06        (o_d_reg[51][6]),
                .reg07        (o_d_reg[51][7]),
                .reg08        (o_d_reg[51][8]),
                .reg09        (o_d_reg[51][9]),
                .reg10        (o_d_reg[51][10]),
                .reg11        (o_d_reg[51][11]),
                .reg12        (o_d_reg[51][12]),
                .reg13        (o_d_reg[51][13]),
                .reg14        (o_d_reg[51][14]),
                .reg15        (o_d_reg[51][15]),
                .reg16        (o_d_reg[51][16]),
                .reg17        (o_d_reg[51][17]),
                .reg18        (o_d_reg[51][18]),
                .reg19        (o_d_reg[51][19]),
                .reg20        (o_d_reg[51][20]),
                .reg21        (o_d_reg[51][21]),
                .reg22        (o_d_reg[51][22]),
                .reg23        (o_d_reg[51][23]),
                .reg24        (o_d_reg[51][24]),
                .reg25        (o_d_reg[51][25]),
                .reg26        (o_d_reg[51][26]),
                .reg27        (o_d_reg[51][27]),
                .reg28        (o_d_reg[51][28]),
                .reg29        (o_d_reg[51][29]),
                .reg30        (o_d_reg[51][30]),
                .reg31        (o_d_reg[51][31]),
                .reg32        (o_d_reg[51][32]),
                .reg33        (o_d_reg[51][33]),
                .reg34        (o_d_reg[51][34]),
                .reg35        (o_d_reg[51][35]),
                .reg36        (o_d_reg[51][36]),
                .reg37        (o_d_reg[51][37]),
                .reg38        (o_d_reg[51][38]),
                .reg39        (o_d_reg[51][39]),
                .reg40        (o_d_reg[51][40]),
                .reg41        (o_d_reg[51][41]),
                .reg42        (o_d_reg[51][42]),
                .reg43        (o_d_reg[51][43]),
                .reg44        (o_d_reg[51][44]),
                .reg45        (o_d_reg[51][45]),
                .reg46        (o_d_reg[51][46]),
                .reg47        (o_d_reg[51][47]),
                .reg48        (o_d_reg[51][48]),
                .reg49        (o_d_reg[51][49]),
                .reg50        (o_d_reg[51][50]),
                .reg51        (o_d_reg[51][51]),
                .reg52        (o_d_reg[51][52])
        );

//last line
regs52
#(
	.DATA_WIDTH(28),
	.REGDEPTH(52)
)
rowBuf52
(
    .clk(clk),
    .rst(rst),
    .din(o_d_rowBuf[REGSNUM-1]),
    .reg43(reg_43_52),
    .reg10(reg_10_52)
);


assign reg_10_01 = o_d_reg[1][10];
assign reg_43_01 = o_d_reg[1][43];
assign reg_12_04 = o_d_reg[4][12];
assign reg_41_04 = o_d_reg[4][41];
assign reg_14_07 = o_d_reg[7][14];
assign reg_39_07 = o_d_reg[7][39];
assign reg_09_09 = o_d_reg[9][9];
assign reg_26_09 = o_d_reg[9][26];
assign reg_27_09 = o_d_reg[9][27];
assign reg_44_09 = o_d_reg[9][44];
assign reg_01_10 = o_d_reg[10][1];
assign reg_16_10 = o_d_reg[10][16];
assign reg_18_10 = o_d_reg[10][18];
assign reg_35_10 = o_d_reg[10][35];
assign reg_37_10 = o_d_reg[10][37];
assign reg_52_10 = o_d_reg[10][52];
assign reg_11_11 = o_d_reg[11][11];
assign reg_26_11 = o_d_reg[11][26];
assign reg_27_11 = o_d_reg[11][27];
assign reg_42_11 = o_d_reg[11][42];
assign reg_04_12 = o_d_reg[12][4] ;
assign reg_19_12 = o_d_reg[12][19];
assign reg_34_12 = o_d_reg[12][34];
assign reg_49_12 = o_d_reg[12][49];
assign reg_13_13 = o_d_reg[13][13];
assign reg_18_13 = o_d_reg[13][18];
assign reg_26_13 = o_d_reg[13][26];
assign reg_27_13 = o_d_reg[13][27];
assign reg_35_13 = o_d_reg[13][35];
assign reg_40_13 = o_d_reg[13][40];
assign reg_07_14 = o_d_reg[14][7] ;
assign reg_20_14 = o_d_reg[14][20];
assign reg_33_14 = o_d_reg[14][33];
assign reg_46_14 = o_d_reg[14][46];
assign reg_15_15 = o_d_reg[15][15];
assign reg_26_15 = o_d_reg[15][26];
assign reg_27_15 = o_d_reg[15][27];
assign reg_38_15 = o_d_reg[15][38];
assign reg_10_16 = o_d_reg[16][10];
assign reg_20_16 = o_d_reg[16][20];
assign reg_21_16 = o_d_reg[16][21];
assign reg_32_16 = o_d_reg[16][32];
assign reg_33_16 = o_d_reg[16][33];
assign reg_43_16 = o_d_reg[16][43];
assign reg_17_17 = o_d_reg[17][17];
assign reg_26_17 = o_d_reg[17][26];
assign reg_27_17 = o_d_reg[17][27];
assign reg_36_17 = o_d_reg[17][36];
assign reg_10_18 = o_d_reg[18][10];
assign reg_13_18 = o_d_reg[18][13];
assign reg_22_18 = o_d_reg[18][22];
assign reg_31_18 = o_d_reg[18][31];
assign reg_40_18 = o_d_reg[18][40];
assign reg_43_18 = o_d_reg[18][43];
assign reg_12_19 = o_d_reg[19][12];
assign reg_19_19 = o_d_reg[19][19];
assign reg_22_19 = o_d_reg[19][22];
assign reg_26_19 = o_d_reg[19][26];
assign reg_27_19 = o_d_reg[19][27];
assign reg_31_19 = o_d_reg[19][31];
assign reg_34_19 = o_d_reg[19][34];
assign reg_41_19 = o_d_reg[19][41];
assign reg_14_20 = o_d_reg[20][14];
assign reg_16_20 = o_d_reg[20][16];
assign reg_23_20 = o_d_reg[20][23];
assign reg_30_20 = o_d_reg[20][30];
assign reg_37_20 = o_d_reg[20][37];
assign reg_39_20 = o_d_reg[20][39];
assign reg_16_21 = o_d_reg[21][16];
assign reg_21_21 = o_d_reg[21][21];
assign reg_26_21 = o_d_reg[21][26];
assign reg_27_21 = o_d_reg[21][27];
assign reg_32_21 = o_d_reg[21][32];
assign reg_37_21 = o_d_reg[21][37];
assign reg_18_22 = o_d_reg[22][18];
assign reg_19_22 = o_d_reg[22][19];
assign reg_24_22 = o_d_reg[22][24];
assign reg_29_22 = o_d_reg[22][29];
assign reg_34_22 = o_d_reg[22][34];
assign reg_35_22 = o_d_reg[22][35];
assign reg_20_23 = o_d_reg[23][20];
assign reg_23_23 = o_d_reg[23][23];
assign reg_26_23 = o_d_reg[23][26];
assign reg_27_23 = o_d_reg[23][27];
assign reg_30_23 = o_d_reg[23][30];
assign reg_33_23 = o_d_reg[23][33];
assign reg_22_24 = o_d_reg[24][22];
assign reg_25_24 = o_d_reg[24][25];
assign reg_28_24 = o_d_reg[24][28];
assign reg_31_24 = o_d_reg[24][31];
assign reg_24_25 = o_d_reg[25][24];
assign reg_29_25 = o_d_reg[25][29];
assign reg_09_26 = o_d_reg[26][9];
assign reg_11_26 = o_d_reg[26][11];
assign reg_13_26 = o_d_reg[26][13];
assign reg_15_26 = o_d_reg[26][15];
assign reg_17_26 = o_d_reg[26][17];
assign reg_19_26 = o_d_reg[26][19];
assign reg_21_26 = o_d_reg[26][21];
assign reg_23_26 = o_d_reg[26][23];
assign reg_26_26 = o_d_reg[26][26];
assign reg_27_26 = o_d_reg[26][27];
assign reg_30_26 = o_d_reg[26][30];
assign reg_32_26 = o_d_reg[26][32];
assign reg_34_26 = o_d_reg[26][34];
assign reg_36_26 = o_d_reg[26][36];
assign reg_38_26 = o_d_reg[26][38];
assign reg_40_26 = o_d_reg[26][40];
assign reg_42_26 = o_d_reg[26][42];
assign reg_44_26 = o_d_reg[26][44];
assign reg_09_27 = o_d_reg[27][9];
assign reg_11_27 = o_d_reg[27][11];
assign reg_13_27 = o_d_reg[27][13];
assign reg_15_27 = o_d_reg[27][15];
assign reg_17_27 = o_d_reg[27][17];
assign reg_19_27 = o_d_reg[27][19];
assign reg_21_27 = o_d_reg[27][21];
assign reg_23_27 = o_d_reg[27][23];
assign reg_26_27 = o_d_reg[27][26];
assign reg_27_27 = o_d_reg[27][27];
assign reg_30_27 = o_d_reg[27][30];
assign reg_32_27 = o_d_reg[27][32];
assign reg_34_27 = o_d_reg[27][34];
assign reg_36_27 = o_d_reg[27][36];
assign reg_38_27 = o_d_reg[27][38];
assign reg_40_27 = o_d_reg[27][40];
assign reg_42_27 = o_d_reg[27][42];
assign reg_44_27 = o_d_reg[27][44];
assign reg_24_28 = o_d_reg[28][24];
assign reg_29_28 = o_d_reg[28][29];
assign reg_22_29 = o_d_reg[29][22];
assign reg_25_29 = o_d_reg[29][25];
assign reg_28_29 = o_d_reg[29][28];
assign reg_31_29 = o_d_reg[29][31];
assign reg_20_30 = o_d_reg[30][20];
assign reg_23_30 = o_d_reg[30][23];
assign reg_26_30 = o_d_reg[30][26];
assign reg_27_30 = o_d_reg[30][27];
assign reg_30_30 = o_d_reg[30][30];
assign reg_33_30 = o_d_reg[30][33];
assign reg_18_31 = o_d_reg[31][18];
assign reg_19_31 = o_d_reg[31][19];
assign reg_24_31 = o_d_reg[31][24];
assign reg_29_31 = o_d_reg[31][29];
assign reg_34_31 = o_d_reg[31][34];
assign reg_35_31 = o_d_reg[31][35];
assign reg_16_32 = o_d_reg[32][16];
assign reg_21_32 = o_d_reg[32][21];
assign reg_26_32 = o_d_reg[32][26];
assign reg_27_32 = o_d_reg[32][27];
assign reg_32_32 = o_d_reg[32][32];
assign reg_37_32 = o_d_reg[32][37];
assign reg_14_33 = o_d_reg[33][14];
assign reg_16_33 = o_d_reg[33][16];
assign reg_23_33 = o_d_reg[33][23];
assign reg_30_33 = o_d_reg[33][30];
assign reg_37_33 = o_d_reg[33][37];
assign reg_39_33 = o_d_reg[33][39];
assign reg_12_34 = o_d_reg[34][12];
assign reg_19_34 = o_d_reg[34][19];
assign reg_22_34 = o_d_reg[34][22];
assign reg_26_34 = o_d_reg[34][26];
assign reg_27_34 = o_d_reg[34][27];
assign reg_31_34 = o_d_reg[34][31];
assign reg_34_34 = o_d_reg[34][34];
assign reg_41_34 = o_d_reg[34][41];
assign reg_10_35 = o_d_reg[35][10];
assign reg_13_35 = o_d_reg[35][13];
assign reg_22_35 = o_d_reg[35][22];
assign reg_31_35 = o_d_reg[35][31];
assign reg_40_35 = o_d_reg[35][40];
assign reg_43_35 = o_d_reg[35][43];
assign reg_17_36 = o_d_reg[36][17];
assign reg_26_36 = o_d_reg[36][26];
assign reg_27_36 = o_d_reg[36][27];
assign reg_36_36 = o_d_reg[36][36];
assign reg_10_37 = o_d_reg[37][10];
assign reg_20_37 = o_d_reg[37][20];
assign reg_21_37 = o_d_reg[37][21];
assign reg_32_37 = o_d_reg[37][32];
assign reg_33_37 = o_d_reg[37][33];
assign reg_43_37 = o_d_reg[37][43];
assign reg_15_38 = o_d_reg[38][15];
assign reg_26_38 = o_d_reg[38][26];
assign reg_27_38 = o_d_reg[38][27];
assign reg_38_38 = o_d_reg[38][38];
assign reg_07_39 = o_d_reg[39][7];
assign reg_20_39 = o_d_reg[39][20];
assign reg_33_39 = o_d_reg[39][33];
assign reg_46_39 = o_d_reg[39][46];
assign reg_13_40 = o_d_reg[40][13];
assign reg_18_40 = o_d_reg[40][18];
assign reg_26_40 = o_d_reg[40][26];
assign reg_27_40 = o_d_reg[40][27];
assign reg_35_40 = o_d_reg[40][35];
assign reg_40_40 = o_d_reg[40][40];
assign reg_04_41 = o_d_reg[41][4];
assign reg_19_41 = o_d_reg[41][19];
assign reg_34_41 = o_d_reg[41][34];
assign reg_49_41 = o_d_reg[41][49];
assign reg_11_42 = o_d_reg[42][11];
assign reg_26_42 = o_d_reg[42][26];
assign reg_27_42 = o_d_reg[42][27];
assign reg_42_42 = o_d_reg[42][42];
assign reg_01_43 = o_d_reg[43][1];
assign reg_16_43 = o_d_reg[43][16];
assign reg_18_43 = o_d_reg[43][18];
assign reg_35_43 = o_d_reg[43][35];
assign reg_37_43 = o_d_reg[43][37];
assign reg_52_43 = o_d_reg[43][52];
assign reg_09_44 = o_d_reg[44][9];
assign reg_26_44 = o_d_reg[44][26];
assign reg_27_44 = o_d_reg[44][27];
assign reg_44_44 = o_d_reg[44][44];
assign reg_14_46 = o_d_reg[46][14];
assign reg_39_46 = o_d_reg[46][39];
assign reg_12_49 = o_d_reg[49][12];
assign reg_41_49 = o_d_reg[49][41];

localparam maxValidLatency = IMAGE_WIDTH*25 + 26;
reg [maxValidLatency-1:0] valid_delay;
integer i;
always @(posedge clk) begin
    for(i=0; i<maxValidLatency-1; i=i+1)
        valid_delay[i+1] <= valid_delay[i];
    valid_delay[0] <= din_valid;
end
assign dout_valid = valid_delay[maxValidLatency-1];

//reg [9:0] delay_col_cnt [maxValidLatency-1:0];
//reg [9:0] delay_row_cnt [maxValidLatency-1:0];
//always @(posedge clk) begin
//    for(i=0; i<maxValidLatency-1; i=i+1)
//        delay_col_cnt[i+1] <= delay_col_cnt[i];
//    delay_col_cnt[0] <= i_col_cnt;
//end
//always @(posedge clk) begin
//    for(i=0; i<maxValidLatency-1; i=i+1)
//        delay_row_cnt[i+1] <= delay_row_cnt[i];
//    delay_row_cnt[0] <= i_row_cnt;
//end

//assign o_col_cnt = delay_col_cnt[maxValidLatency-1];
//assign o_row_cnt = delay_row_cnt[maxValidLatency-1];


endmodule
